CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 23 100 9
38 96 1497 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 96 1497 799
143654930 0
0
6 Title:
5 Name:
0
0
0
29
13 Logic Switch~
5 945 47 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 946 92 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 946 136 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -18 8 -10
2 A3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 946 180 0 1 11
0 21
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 1180 170 0 1 11
0 22
0
0 0 21360 512
2 0V
-7 -16 7 -8
2 B1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 1181 123 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 B2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 1181 81 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 B3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 1181 43 0 1 11
0 25
0
0 0 21360 512
2 0V
-7 -16 7 -8
2 B4
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3747 0 0
0
0
13 Logic Switch~
5 1349 107 0 1 11
0 5
0
0 0 21360 512
2 0V
-8 -17 6 -9
1 M
-4 -26 3 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3549 0 0
0
0
12 2-Input XOR~
16 1021 557 0 3 22
0 6 5 4
0
0 0 624 512
6 74LS86
-21 -24 21 -16
3 U8A
0 -25 21 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -1493283793
65 0 0 0 4 1 5 0
1 U
7931 0 0
0
0
11 2-Input OR~
1 1068 551 0 3 22
0 8 7 6
0
0 0 880 512
6 74LS32
-9 -25 33 -17
3 U4B
1 -35 22 -27
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 -1493283793
65 0 0 0 4 2 3 0
1 U
9325 0 0
0
0
7 Ground~
168 429 326 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8903 0 0
0
0
12 2-Input AND~
0 1160 502 0 3 22
0 14 13 7
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U7A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -1224782786
65 0 0 0 4 1 4 0
1 U
3834 0 0
0
0
11 2-Input OR~
1 1160 416 0 3 22
0 15 16 14
0
0 0 880 270
6 74LS32
29 -2 71 6
3 U4A
39 -12 60 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -1375843292
65 0 0 0 4 1 3 0
1 U
3363 0 0
0
0
7 Ground~
168 951 447 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7668 0 0
0
0
6 74LS83
105 896 372 0 14 29
0 13 16 15 17 2 4 4 2 2
12 11 10 9 46
0
0 0 13040 512
7 74LS83A
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
4718 0 0
0
0
6 74LS83
105 1035 245 0 14 29
0 21 20 19 18 26 27 28 29 5
13 16 15 17 8
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
2 U6
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3874 0 0
0
0
12 2-Input XOR~
16 1150 176 0 3 22
0 5 22 29
0
0 0 624 180
6 74LS86
-21 -24 21 -16
3 U5D
0 -25 21 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 2 0
1 U
6671 0 0
0
0
12 2-Input XOR~
16 1149 130 0 3 22
0 23 5 28
0
0 0 624 512
6 74LS86
-21 -24 21 -16
3 U5C
0 -25 21 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 2 0
1 U
3789 0 0
0
0
12 2-Input XOR~
16 1149 87 0 3 22
0 5 24 27
0
0 0 624 180
6 74LS86
-21 -24 21 -16
3 U5B
0 -25 21 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 2 0
1 U
4871 0 0
0
0
12 2-Input XOR~
16 1150 49 0 3 22
0 5 25 26
0
0 0 624 180
6 74LS86
-21 -24 21 -16
3 U5A
0 -25 21 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 2 0
1 U
3750 0 0
0
0
9 CA 7-Seg~
184 540 181 0 18 19
10 36 35 34 33 32 31 30 47 37
0 0 2 0 0 2 0 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
8778 0 0
0
0
2 +V
167 540 77 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
538 0 0
0
0
6 74LS47
187 525 262 0 14 29
0 12 11 10 9 48 49 30 31 32
33 34 35 36 50
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U2
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
6843 0 0
0
0
6 74LS47
187 389 262 0 14 29
0 2 2 2 4 51 52 38 39 40
41 42 43 44 53
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U1
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3136 0 0
0
0
2 +V
167 404 77 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5950 0 0
0
0
9 CA 7-Seg~
184 404 181 0 18 19
10 44 43 42 41 40 39 38 54 45
2 0 0 2 2 2 2 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
5670 0 0
0
0
9 Resistor~
219 540 115 0 4 5
0 37 3 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6828 0 0
0
0
9 Resistor~
219 404 115 0 4 5
0 45 3 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6735 0 0
0
0
60
4 3 4 0 0 8320 0 25 10 0 0 3
403 299
403 557
994 557
0 3 4 0 0 0 0 0 10 7 0 4
928 386
998 386
998 557
994 557
1 2 5 0 0 4224 0 9 10 0 0 3
1337 107
1337 563
1042 563
1 3 6 0 0 4224 0 10 11 0 0 2
1042 551
1041 551
3 2 7 0 0 8320 0 13 11 0 0 3
1158 525
1158 557
1086 557
14 1 8 0 0 4224 0 17 11 0 0 5
1078 279
1078 532
1109 532
1109 545
1086 545
7 6 4 0 0 0 0 16 16 0 0 2
928 390
928 381
4 13 9 0 0 8320 0 24 16 0 0 3
539 299
539 390
864 390
3 12 10 0 0 8320 0 24 16 0 0 3
548 299
548 381
864 381
2 11 11 0 0 8320 0 24 16 0 0 3
557 299
557 372
864 372
1 10 12 0 0 8320 0 24 16 0 0 3
566 299
566 363
864 363
1 1 2 0 0 4096 0 25 12 0 0 4
430 299
430 312
429 312
429 320
2 1 2 0 0 0 0 25 25 0 0 2
421 299
430 299
3 2 2 0 0 0 0 25 25 0 0 2
412 299
421 299
10 2 13 0 0 4224 0 17 13 0 0 4
1024 279
1024 472
1152 472
1152 480
3 1 14 0 0 4224 0 14 13 0 0 4
1163 446
1163 472
1164 472
1164 480
12 1 15 0 0 8320 0 17 14 0 0 4
1042 279
1042 386
1169 386
1169 401
11 2 16 0 0 8320 0 17 14 0 0 4
1033 279
1033 386
1157 386
1157 401
8 1 2 0 0 8192 0 16 15 0 0 3
928 399
951 399
951 441
5 1 2 0 0 8320 0 16 15 0 0 3
928 372
951 372
951 441
9 1 2 0 0 0 0 16 15 0 0 3
928 417
951 417
951 441
13 4 17 0 0 8320 0 17 16 0 0 3
1051 279
1051 363
928 363
12 3 15 0 0 0 0 17 16 0 0 3
1042 279
1042 354
928 354
11 2 16 0 0 0 0 17 16 0 0 3
1033 279
1033 345
928 345
10 1 13 0 0 0 0 17 16 0 0 3
1024 279
1024 336
928 336
1 4 18 0 0 8320 0 1 17 0 0 3
957 47
1024 47
1024 215
1 3 19 0 0 8320 0 2 17 0 0 3
958 92
1015 92
1015 215
1 2 20 0 0 8320 0 3 17 0 0 3
958 136
1006 136
1006 215
1 1 21 0 0 4224 0 4 17 0 0 3
958 180
997 180
997 215
9 1 5 0 0 0 0 17 9 0 0 3
1078 215
1078 107
1337 107
1 1 5 0 0 0 0 18 9 0 0 4
1171 182
1331 182
1331 107
1337 107
2 0 5 0 0 0 0 19 0 0 34 4
1170 136
1326 136
1326 105
1331 105
1 0 5 0 0 0 0 20 0 0 34 2
1170 93
1331 93
1 1 5 0 0 0 0 21 9 0 0 4
1171 55
1331 55
1331 107
1337 107
1 2 22 0 0 4224 0 5 18 0 0 2
1168 170
1171 170
1 1 23 0 0 4224 0 6 19 0 0 3
1169 123
1169 124
1170 124
1 2 24 0 0 4224 0 7 20 0 0 2
1169 81
1170 81
1 2 25 0 0 4224 0 8 21 0 0 2
1169 43
1171 43
3 5 26 0 0 8320 0 21 17 0 0 3
1123 49
1033 49
1033 215
3 6 27 0 0 8320 0 20 17 0 0 3
1122 87
1042 87
1042 215
3 7 28 0 0 8320 0 19 17 0 0 3
1122 130
1051 130
1051 215
3 8 29 0 0 4224 0 18 17 0 0 3
1123 176
1060 176
1060 215
7 7 30 0 0 8320 0 24 22 0 0 4
566 229
566 225
555 225
555 217
8 6 31 0 0 8320 0 24 22 0 0 4
557 229
557 225
549 225
549 217
9 5 32 0 0 12416 0 24 22 0 0 4
548 229
548 225
543 225
543 217
10 4 33 0 0 12416 0 24 22 0 0 4
539 229
539 225
537 225
537 217
11 3 34 0 0 12416 0 24 22 0 0 4
530 229
530 225
531 225
531 217
12 2 35 0 0 12416 0 24 22 0 0 4
521 229
521 225
525 225
525 217
13 1 36 0 0 12416 0 24 22 0 0 4
512 229
512 225
519 225
519 217
1 2 3 0 0 4224 0 23 28 0 0 2
540 86
540 97
1 9 37 0 0 4224 0 28 22 0 0 2
540 133
540 145
7 7 38 0 0 8320 0 25 27 0 0 4
430 229
430 225
419 225
419 217
8 6 39 0 0 8320 0 25 27 0 0 4
421 229
421 225
413 225
413 217
9 5 40 0 0 12416 0 25 27 0 0 4
412 229
412 225
407 225
407 217
10 4 41 0 0 12416 0 25 27 0 0 4
403 229
403 225
401 225
401 217
11 3 42 0 0 12416 0 25 27 0 0 4
394 229
394 225
395 225
395 217
12 2 43 0 0 12416 0 25 27 0 0 4
385 229
385 225
389 225
389 217
13 1 44 0 0 12416 0 25 27 0 0 4
376 229
376 225
383 225
383 217
1 2 3 0 0 0 0 26 29 0 0 2
404 86
404 97
1 9 45 0 0 4224 0 29 27 0 0 2
404 133
404 145
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
