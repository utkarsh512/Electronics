CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 130 9
38 96 1497 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 96 1497 799
143654930 0
0
6 Title:
5 Name:
0
0
0
28
7 Ground~
168 183 208 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 512 0 0 0 0
3 GND
8953 0 0
0
0
11 2-Input OR~
1 457 453 0 3 22
0 5 6 4
0
0 0 880 512
6 74LS32
-9 -25 33 -17
3 U8C
1 -35 22 -27
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 912162011
65 0 0 0 4 3 4 0
1 U
4441 0 0
0
0
11 4-Input OR~
219 455 355 0 5 12
0 8 5 9 10 7
0
0 0 624 512
4 4072
-14 -24 14 -16
3 U7B
1 -25 22 -17
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 912162011
65 0 0 0 2 2 3 0
1 U
3618 0 0
0
0
11 3-Input OR~
86 454 273 0 4 22
0 8 12 10 11
0
0 0 624 512
4 4075
-14 -28 14 -20
3 U9C
1 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 11 12 13 10 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 3 5 0
1 U
6153 0 0
0
0
11 3-Input OR~
86 451 201 0 4 22
0 9 10 14 13
0
0 0 624 512
4 4075
-14 -28 14 -20
3 U9B
1 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 8 9 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 2 5 0
1 U
5394 0 0
0
0
7 Ground~
168 215 432 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7734 0 0
0
0
11 2-Input OR~
1 370 397 0 3 22
0 6 5 15
0
0 0 880 180
6 74LS32
-9 -25 33 -17
3 U8B
1 -35 22 -27
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 912162011
65 0 0 0 4 2 4 0
1 U
9914 0 0
0
0
11 3-Input OR~
86 368 316 0 4 22
0 5 9 10 16
0
0 0 624 512
4 4075
-14 -28 14 -20
3 U9A
1 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 3 5 6 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 5 0
1 U
3747 0 0
0
0
11 2-Input OR~
1 366 239 0 3 22
0 10 12 17
0
0 0 880 180
6 74LS32
-9 -25 33 -17
3 U8A
1 -35 22 -27
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 593460431
65 0 0 0 4 1 4 0
1 U
3549 0 0
0
0
11 4-Input OR~
219 365 163 0 5 12
0 14 10 9 8 18
0
0 0 624 180
4 4072
-14 -24 14 -16
3 U7A
1 -25 22 -17
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 643792074
65 0 0 0 2 1 3 0
1 U
7931 0 0
0
0
7 74LS157
122 183 310 0 14 29
0 43 18 13 17 11 16 7 15 4
2 22 21 20 19
0
0 0 13040 512
7 74LS157
-24 -60 25 -52
2 U6
-13 -61 1 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 512 1 0 0 0
1 U
9325 0 0
0
0
6 74LS47
187 81 230 0 14 29
0 22 21 20 19 44 45 23 24 25
26 27 28 29 46
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U1
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
8903 0 0
0
0
2 +V
167 96 45 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3834 0 0
0
0
9 CA 7-Seg~
184 96 149 0 18 19
10 29 28 27 26 25 24 23 47 30
2 2 2 0 0 2 0 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3363 0 0
0
0
9 Inverter~
13 635 477 0 2 22
0 38 6
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U5B
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
7668 0 0
0
0
9 Inverter~
13 636 449 0 2 22
0 37 14
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U5A
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
4718 0 0
0
0
9 Inverter~
13 636 426 0 2 22
0 36 10
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U4F
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
3874 0 0
0
0
9 Inverter~
13 636 402 0 2 22
0 35 9
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U4E
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
6671 0 0
0
0
9 Inverter~
13 635 377 0 2 22
0 34 5
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U4D
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
3789 0 0
0
0
9 Inverter~
13 635 352 0 2 22
0 33 48
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U4C
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 512 6 3 1 0
1 U
4871 0 0
0
0
9 Inverter~
13 635 324 0 2 22
0 32 12
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U4B
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3750 0 0
0
0
9 Inverter~
13 635 298 0 2 22
0 31 8
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U4A
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
8778 0 0
0
0
7 Ground~
168 855 205 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
538 0 0
0
0
7 74LS138
19 778 252 0 14 29
0 41 40 39 49 2 2 31 32 33
34 35 36 37 38
0
0 0 13296 782
7 74LS138
50 -2 99 6
2 U3
68 -12 82 -4
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 512 1 0 0 0
1 U
6843 0 0
0
0
7 Pulser~
4 823 95 0 10 12
0 50 51 42 52 0 0 5 5 4
7
0
0 0 4656 512
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3136 0 0
0
0
7 Ground~
168 707 115 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5950 0 0
0
0
6 74LS93
109 756 157 0 8 17
0 2 2 42 39 53 41 40 39
0
0 0 13040 782
6 74LS93
-21 -35 21 -27
2 U2
28 0 42 8
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 512 1 0 0 0
1 U
5670 0 0
0
0
9 Resistor~
219 96 83 0 4 5
0 30 3 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6828 0 0
0
0
62
3 9 4 0 0 4224 0 2 11 0 0 4
430 453
229 453
229 346
209 346
1 2 5 0 0 4096 0 2 19 0 0 4
475 447
612 447
612 377
620 377
2 2 6 0 0 4096 0 2 15 0 0 4
475 459
612 459
612 477
620 477
5 7 7 0 0 4224 0 3 11 0 0 4
428 355
223 355
223 328
209 328
2 1 8 0 0 4096 0 22 3 0 0 4
620 298
496 298
496 346
474 346
2 2 5 0 0 0 0 19 3 0 0 4
620 377
496 377
496 352
473 352
2 3 9 0 0 4096 0 18 3 0 0 4
621 402
496 402
496 358
473 358
2 4 10 0 0 4096 0 17 3 0 0 4
621 426
496 426
496 364
474 364
4 5 11 0 0 4224 0 4 11 0 0 4
427 273
223 273
223 310
209 310
1 2 8 0 0 4096 0 4 22 0 0 4
473 264
612 264
612 298
620 298
2 2 12 0 0 4096 0 4 21 0 0 4
472 273
612 273
612 324
620 324
2 3 10 0 0 8192 0 17 4 0 0 4
621 426
495 426
495 282
473 282
4 3 13 0 0 4224 0 5 11 0 0 4
424 201
223 201
223 292
209 292
1 2 9 0 0 8192 0 5 18 0 0 4
470 192
613 192
613 402
621 402
2 2 10 0 0 8192 0 5 17 0 0 4
469 201
613 201
613 426
621 426
3 2 14 0 0 8192 0 5 16 0 0 4
470 210
613 210
613 449
621 449
10 1 2 0 0 8320 0 11 6 0 0 5
215 355
219 355
219 418
215 418
215 426
3 8 15 0 0 4224 0 7 11 0 0 4
343 397
223 397
223 337
209 337
2 2 5 0 0 4096 0 7 19 0 0 4
388 391
612 391
612 377
620 377
1 2 6 0 0 4224 0 7 15 0 0 4
388 403
612 403
612 477
620 477
4 6 16 0 0 4224 0 8 11 0 0 4
341 316
223 316
223 319
209 319
1 2 5 0 0 4224 0 8 19 0 0 4
387 307
612 307
612 377
620 377
2 2 9 0 0 4096 0 8 18 0 0 4
386 316
613 316
613 402
621 402
3 2 10 0 0 4096 0 8 17 0 0 4
387 325
613 325
613 426
621 426
3 4 17 0 0 4224 0 9 11 0 0 4
339 239
223 239
223 301
209 301
2 2 12 0 0 4224 0 21 9 0 0 4
620 324
406 324
406 233
384 233
2 1 10 0 0 0 0 17 9 0 0 4
621 426
406 426
406 245
384 245
4 2 8 0 0 4224 0 10 22 0 0 4
384 154
612 154
612 298
620 298
3 2 9 0 0 8320 0 10 18 0 0 4
383 160
613 160
613 402
621 402
2 2 10 0 0 8320 0 10 17 0 0 4
383 166
613 166
613 426
621 426
1 2 14 0 0 8320 0 10 16 0 0 4
384 172
613 172
613 449
621 449
5 2 18 0 0 8320 0 10 11 0 0 4
338 163
223 163
223 283
209 283
4 14 19 0 0 4224 0 12 11 0 0 3
95 267
95 346
145 346
3 13 20 0 0 4224 0 12 11 0 0 3
104 267
104 328
145 328
2 12 21 0 0 4224 0 12 11 0 0 3
113 267
113 310
145 310
1 11 22 0 0 4224 0 12 11 0 0 3
122 267
122 292
145 292
7 7 23 0 0 8336 0 12 14 0 0 4
122 197
122 193
111 193
111 185
8 6 24 0 0 8336 0 12 14 0 0 4
113 197
113 193
105 193
105 185
9 5 25 0 0 12432 0 12 14 0 0 4
104 197
104 193
99 193
99 185
10 4 26 0 0 12432 0 12 14 0 0 4
95 197
95 193
93 193
93 185
11 3 27 0 0 12432 0 12 14 0 0 4
86 197
86 193
87 193
87 185
12 2 28 0 0 12432 0 12 14 0 0 4
77 197
77 193
81 193
81 185
13 1 29 0 0 12432 0 12 14 0 0 4
68 197
68 193
75 193
75 185
1 2 3 0 0 4240 0 13 28 0 0 2
96 54
96 65
1 9 30 0 0 4240 0 28 14 0 0 2
96 101
96 113
7 1 31 0 0 8320 0 24 22 0 0 3
753 288
753 298
656 298
8 1 32 0 0 8320 0 24 21 0 0 3
762 288
762 324
656 324
9 1 33 0 0 8320 0 24 20 0 0 3
771 288
771 352
656 352
10 1 34 0 0 8320 0 24 19 0 0 3
780 288
780 377
656 377
11 1 35 0 0 8320 0 24 18 0 0 3
789 288
789 402
657 402
12 1 36 0 0 8320 0 24 17 0 0 3
798 288
798 426
657 426
13 1 37 0 0 4224 0 24 16 0 0 3
807 288
807 449
657 449
14 1 38 0 0 4224 0 24 15 0 0 3
816 288
816 477
656 477
6 1 2 0 0 0 0 24 23 0 0 4
816 212
816 191
855 191
855 199
5 1 2 0 0 128 0 24 23 0 0 4
807 212
807 191
855 191
855 199
8 4 39 0 0 12416 0 27 27 0 0 6
770 193
770 197
785 197
785 115
770 115
770 123
8 3 39 0 0 0 0 27 24 0 0 4
770 193
770 203
771 203
771 218
7 2 40 0 0 12416 0 27 24 0 0 4
761 193
761 203
762 203
762 218
6 1 41 0 0 12416 0 27 24 0 0 4
752 193
752 203
753 203
753 218
3 3 42 0 0 8320 0 27 25 0 0 3
761 123
761 86
799 86
0 1 2 0 0 0 0 0 26 62 0 4
747 129
747 85
707 85
707 109
1 2 2 0 0 0 0 27 27 0 0 2
743 129
752 129
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
285 18 405 42
293 25 405 41
14 18EC30048 & 46
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
