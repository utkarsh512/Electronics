CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
38 96 1497 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 96 1497 799
143654930 0
0
6 Title:
5 Name:
0
0
0
41
13 Logic Switch~
5 646 44 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-6 -16 8 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 639 263 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-6 -16 8 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 670 340 0 1 11
0 6
0
0 0 21360 512
2 0V
-15 -11 -1 -3
2 V9
-14 -20 0 -12
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 659 306 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-6 -16 8 -8
2 V8
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 695 363 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
16 -19 30 -11
2 V7
15 -27 29 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 696 400 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-6 -16 8 -8
2 V3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 697 441 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-6 -16 8 -8
2 V2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 700 489 0 10 11
0 27 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-6 -16 8 -8
2 V1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3747 0 0
0
0
13 Logic Switch~
5 326 472 0 1 11
0 50
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3549 0 0
0
0
13 Logic Switch~
5 175 423 0 10 11
0 48 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7931 0 0
0
0
14 Logic Display~
6 528 226 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9325 0 0
0
0
14 Logic Display~
6 446 281 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8903 0 0
0
0
14 Logic Display~
6 468 282 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3834 0 0
0
0
14 Logic Display~
6 490 284 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3363 0 0
0
0
14 Logic Display~
6 512 286 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7668 0 0
0
0
14 Logic Display~
6 264 98 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4718 0 0
0
0
14 Logic Display~
6 294 99 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3874 0 0
0
0
14 Logic Display~
6 327 100 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6671 0 0
0
0
14 Logic Display~
6 359 101 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3789 0 0
0
0
14 Logic Display~
6 390 102 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4871 0 0
0
0
14 Logic Display~
6 420 103 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3750 0 0
0
0
14 Logic Display~
6 451 104 0 1 2
10 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8778 0 0
0
0
8 2-In OR~
219 465 452 0 3 22
0 21 22 23
0
0 0 624 90
6 74LS32
-21 -24 21 -16
3 U6D
28 -3 49 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 -1281517838
65 0 0 0 4 4 2 0
1 U
538 0 0
0
0
8 2-In OR~
219 517 527 0 3 22
0 10 9 21
0
0 0 624 180
6 74LS32
-21 -24 21 -16
3 U6C
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 2 0
1 U
6843 0 0
0
0
8 2-In OR~
219 517 485 0 3 22
0 8 7 22
0
0 0 624 180
6 74LS32
-21 -24 21 -16
3 U6B
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 -1281517838
65 0 0 0 4 2 2 0
1 U
3136 0 0
0
0
9 2-In AND~
219 505 377 0 3 22
0 20 23 5
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 -1080191234
65 0 0 0 4 2 3 0
1 U
5950 0 0
0
0
7 74LS193
137 593 395 0 14 29
0 4 5 11 6 24 25 26 27 51
52 7 8 9 10
0
0 0 13040 512
7 74LS193
-24 -51 25 -43
2 U8
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
5670 0 0
0
0
7 Ground~
168 850 138 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6828 0 0
0
0
7 74LS273
150 604 159 0 18 37
0 3 5 28 29 30 31 32 33 34
35 12 13 14 15 16 17 18 19
0
0 0 13040 512
7 74LS273
-24 -60 25 -52
2 U5
-13 -61 1 -53
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
6735 0 0
0
0
7 Ground~
168 814 271 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8365 0 0
0
0
6 74LS83
105 766 215 0 14 29
0 16 17 18 19 37 38 39 40 2
32 33 34 35 36
0
0 0 13040 512
7 74LS83A
-24 -60 25 -52
2 U4
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
4132 0 0
0
0
6 74LS83
105 765 84 0 14 29
0 12 13 14 15 2 2 2 2 36
28 29 30 31 53
0
0 0 13040 512
7 74LS83A
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
4551 0 0
0
0
7 Ground~
168 921 26 0 1 3
0 2
0
0 0 53360 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3635 0 0
0
0
7 Ground~
168 1032 29 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3973 0 0
0
0
7 74LS173
129 982 207 0 14 29
0 2 2 2 45 41 42 43 44 2
2 37 38 39 40
0
0 0 13040 512
7 74LS173
-24 -51 25 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
3851 0 0
0
0
14 Logic Display~
6 482 106 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8383 0 0
0
0
7 Pulser~
4 159 311 0 10 12
0 54 55 47 56 0 0 5 5 3
8
0
0 0 4656 0
0
2 V6
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9334 0 0
0
0
9 2-In AND~
219 323 355 0 3 22
0 47 48 49
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 2065446846
65 0 0 0 4 1 3 0
1 U
7471 0 0
0
0
8 2-In OR~
219 423 368 0 3 22
0 49 50 20
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U6A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 1746679725
65 0 0 0 4 1 2 0
1 U
3334 0 0
0
0
7 Buffer~
58 1082 207 0 2 22
0 46 45
0
0 0 624 180
4 4050
-14 -19 14 -11
3 U1A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 1 0
1 U
3559 0 0
0
0
10 Ascii Key~
169 1211 217 0 11 12
0 44 43 42 41 57 58 59 46 0
0 58
0
0 0 4656 270
0
4 KBD1
-12 -38 16 -30
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
984 0 0
0
0
72
1 1 3 0 0 8320 0 29 1 0 0 6
636 123
640 123
640 54
631 54
631 44
634 44
1 1 4 0 0 8320 0 27 2 0 0 6
625 368
635 368
635 273
624 273
624 263
627 263
1 3 5 0 0 4096 0 11 26 0 0 5
528 244
528 358
534 358
534 377
526 377
4 1 6 0 0 8320 0 27 3 0 0 4
625 395
652 395
652 340
658 340
1 11 7 0 0 8320 0 12 27 0 0 5
446 299
446 327
539 327
539 404
561 404
1 12 8 0 0 8320 0 13 27 0 0 4
468 300
468 320
561 320
561 413
1 13 9 0 0 12416 0 14 27 0 0 5
490 302
490 314
543 314
543 422
561 422
1 14 10 0 0 12416 0 15 27 0 0 5
512 304
512 309
547 309
547 431
561 431
3 1 11 0 0 8320 0 27 4 0 0 4
631 386
641 386
641 306
647 306
1 11 12 0 0 8320 0 16 29 0 0 3
264 116
264 141
566 141
1 12 13 0 0 8320 0 17 29 0 0 3
294 117
294 150
566 150
1 13 14 0 0 8192 0 18 29 0 0 3
327 118
327 159
566 159
1 14 15 0 0 8192 0 19 29 0 0 3
359 119
359 168
566 168
1 15 16 0 0 8192 0 20 29 0 0 3
390 120
390 177
566 177
1 16 17 0 0 8192 0 21 29 0 0 3
420 121
420 186
566 186
1 17 18 0 0 8192 0 22 29 0 0 3
451 122
451 195
566 195
1 18 19 0 0 8192 0 36 29 0 0 3
482 124
482 204
566 204
3 2 5 0 0 8320 0 26 29 0 0 6
526 377
551 377
551 103
644 103
644 132
630 132
3 2 5 0 0 0 0 26 27 0 0 6
526 377
551 377
551 348
639 348
639 377
625 377
3 1 20 0 0 4224 0 39 26 0 0 2
456 368
481 368
1 3 21 0 0 4224 0 23 24 0 0 3
459 468
459 527
490 527
2 3 22 0 0 4224 0 23 25 0 0 3
477 468
477 485
490 485
3 2 23 0 0 4224 0 23 26 0 0 3
468 422
468 386
481 386
14 1 10 0 0 0 0 27 24 0 0 6
561 431
551 431
551 466
555 466
555 536
536 536
13 2 9 0 0 0 0 27 24 0 0 6
561 422
551 422
551 466
555 466
555 518
536 518
12 1 8 0 0 0 0 27 25 0 0 6
561 413
551 413
551 466
555 466
555 494
536 494
11 2 7 0 0 0 0 27 25 0 0 6
561 404
551 404
551 466
555 466
555 476
536 476
5 1 24 0 0 4224 0 27 5 0 0 4
625 404
677 404
677 363
683 363
6 1 25 0 0 4224 0 27 6 0 0 4
625 413
678 413
678 400
684 400
7 1 26 0 0 4224 0 27 7 0 0 4
625 422
679 422
679 441
685 441
8 1 27 0 0 8320 0 27 8 0 0 4
625 431
682 431
682 489
688 489
18 4 19 0 0 8320 0 29 31 0 0 3
566 204
566 206
798 206
17 3 18 0 0 8320 0 29 31 0 0 3
566 195
566 197
798 197
16 2 17 0 0 8320 0 29 31 0 0 3
566 186
566 188
798 188
15 1 16 0 0 8320 0 29 31 0 0 3
566 177
566 179
798 179
14 4 15 0 0 12416 0 29 32 0 0 6
566 168
562 168
562 28
805 28
805 75
797 75
13 3 14 0 0 12416 0 29 32 0 0 6
566 159
562 159
562 28
805 28
805 66
797 66
12 2 13 0 0 0 0 29 32 0 0 6
566 150
562 150
562 28
805 28
805 57
797 57
11 1 12 0 0 0 0 29 32 0 0 6
566 141
562 141
562 28
805 28
805 48
797 48
5 1 2 0 0 4096 0 32 28 0 0 3
797 84
850 84
850 132
6 1 2 0 0 0 0 32 28 0 0 3
797 93
850 93
850 132
7 1 2 0 0 0 0 32 28 0 0 3
797 102
850 102
850 132
8 1 2 0 0 0 0 32 28 0 0 3
797 111
850 111
850 132
10 3 28 0 0 4224 0 32 29 0 0 4
733 75
644 75
644 141
630 141
11 4 29 0 0 4224 0 32 29 0 0 4
733 84
644 84
644 150
630 150
12 5 30 0 0 4224 0 32 29 0 0 4
733 93
644 93
644 159
630 159
13 6 31 0 0 4224 0 32 29 0 0 4
733 102
644 102
644 168
630 168
10 7 32 0 0 4224 0 31 29 0 0 4
734 206
644 206
644 177
630 177
11 8 33 0 0 4224 0 31 29 0 0 4
734 215
644 215
644 186
630 186
12 9 34 0 0 4224 0 31 29 0 0 4
734 224
644 224
644 195
630 195
13 10 35 0 0 4224 0 31 29 0 0 4
734 233
644 233
644 204
630 204
14 9 36 0 0 8320 0 31 32 0 0 6
734 260
729 260
729 28
805 28
805 129
797 129
9 1 2 0 0 0 0 31 30 0 0 3
798 260
814 260
814 265
11 5 37 0 0 4224 0 35 31 0 0 4
950 216
806 216
806 215
798 215
12 6 38 0 0 4224 0 35 31 0 0 4
950 225
806 225
806 224
798 224
13 7 39 0 0 4224 0 35 31 0 0 4
950 234
806 234
806 233
798 233
14 8 40 0 0 4224 0 35 31 0 0 4
950 243
806 243
806 242
798 242
10 1 2 0 0 8192 0 35 33 0 0 3
944 189
921 189
921 34
9 1 2 0 0 0 0 35 33 0 0 3
944 180
921 180
921 34
3 1 2 0 0 8320 0 35 34 0 0 3
1020 198
1032 198
1032 37
2 1 2 0 0 0 0 35 34 0 0 3
1020 189
1032 189
1032 37
1 1 2 0 0 0 0 35 34 0 0 3
1014 180
1032 180
1032 37
4 5 41 0 0 4224 0 41 35 0 0 4
1187 220
1024 220
1024 216
1014 216
3 6 42 0 0 4224 0 41 35 0 0 4
1187 226
1024 226
1024 225
1014 225
2 7 43 0 0 4224 0 41 35 0 0 4
1187 232
1024 232
1024 234
1014 234
1 8 44 0 0 4224 0 41 35 0 0 4
1187 238
1024 238
1024 243
1014 243
4 2 45 0 0 4224 0 35 40 0 0 2
1014 207
1067 207
1 8 46 0 0 12416 0 40 41 0 0 4
1097 207
1109 207
1109 196
1187 196
3 1 47 0 0 4224 0 37 38 0 0 4
183 302
291 302
291 346
299 346
1 2 48 0 0 4224 0 10 38 0 0 4
187 423
291 423
291 364
299 364
3 1 49 0 0 4224 0 38 39 0 0 4
344 355
402 355
402 359
410 359
1 2 50 0 0 8320 0 9 39 0 0 4
338 472
402 472
402 377
410 377
10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
674 322 698 346
684 330 700 346
2 MR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
661 288 741 312
671 296 743 312
9 PL-ENABLE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
433 231 505 255
443 239 507 255
8 DEBUGGER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
716 406 804 430
726 414 806 430
10 MULTIPLIER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
1164 129 1268 153
1174 137 1270 153
12 MULTIPLICAND
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
335 48 399 72
345 56 401 72
7 PRODUCT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
131 452 219 476
141 460 221 476
10 AUTO-CLOCK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
271 499 375 523
281 507 377 523
12 MANUAL CLOCK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
150 433 182 457
160 441 184 457
3 SW2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
301 477 333 501
311 485 335 501
3 SW3
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
