CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 40 23 130 9
38 96 1497 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 96 1497 799
143654930 0
0
6 Title:
5 Name:
0
0
0
26
7 Pulser~
4 837 488 0 10 12
0 56 57 4 58 0 0 5 5 6
7
0
0 0 4656 0
0
2 V5
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
8953 0 0
0
0
7 Ground~
168 349 303 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4441 0 0
0
0
7 Ground~
168 903 420 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3618 0 0
0
0
6 74LS90
107 896 365 0 10 21
0 2 2 2 2 4 11 5 12 13
11
0
0 0 13040 602
6 74LS90
-21 -51 21 -43
2 U8
40 -11 54 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
6153 0 0
0
0
6 74LS47
187 860 264 0 14 29
0 5 12 13 11 59 8 14 15 16
17 18 19 20 60
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U7
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
5394 0 0
0
0
2 +V
167 875 79 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V4
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7734 0 0
0
0
9 CA 7-Seg~
184 875 183 0 18 19
10 20 19 18 17 16 15 14 61 21
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP4
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
9914 0 0
0
0
7 Ground~
168 740 421 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3747 0 0
0
0
6 74LS90
107 733 366 0 10 21
0 2 2 2 2 5 22 6 23 24
22
0
0 0 13040 602
6 74LS90
-21 -51 21 -43
2 U6
40 -11 54 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
3549 0 0
0
0
6 74LS47
187 697 265 0 14 29
0 6 23 24 22 62 9 25 26 27
28 29 30 31 8
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U5
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
7931 0 0
0
0
2 +V
167 712 80 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9325 0 0
0
0
9 CA 7-Seg~
184 712 184 0 18 19
10 31 30 29 28 27 26 25 63 32
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP3
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
8903 0 0
0
0
7 Ground~
168 432 418 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3834 0 0
0
0
6 74LS90
107 425 363 0 10 21
0 2 2 2 2 7 33 35 34 36
33
0
0 0 13040 602
6 74LS90
-21 -51 21 -43
2 U3
40 -11 54 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
3363 0 0
0
0
6 74LS47
187 389 262 0 14 29
0 35 34 36 33 64 2 37 38 39
40 41 42 43 10
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U1
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
7668 0 0
0
0
2 +V
167 404 77 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4718 0 0
0
0
9 CA 7-Seg~
184 404 181 0 18 19
10 43 42 41 40 39 38 37 65 44
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3874 0 0
0
0
9 CA 7-Seg~
184 552 185 0 18 19
10 54 53 52 51 50 49 48 66 55
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
6671 0 0
0
0
2 +V
167 552 81 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3789 0 0
0
0
6 74LS47
187 537 266 0 14 29
0 7 46 47 45 67 10 48 49 50
51 52 53 54 9
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U4
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
4871 0 0
0
0
6 74LS90
107 573 367 0 10 21
0 2 2 2 2 6 45 7 46 47
45
0
0 0 13040 602
6 74LS90
-21 -51 21 -43
2 U2
40 -11 54 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
3750 0 0
0
0
7 Ground~
168 580 422 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8778 0 0
0
0
9 Resistor~
219 875 117 0 4 5
0 21 3 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
538 0 0
0
0
9 Resistor~
219 712 118 0 4 5
0 32 3 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6843 0 0
0
0
9 Resistor~
219 404 115 0 4 5
0 44 3 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3136 0 0
0
0
9 Resistor~
219 552 119 0 4 5
0 55 3 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5950 0 0
0
0
80
5 3 4 0 0 4224 0 4 1 0 0 3
872 397
872 479
861 479
5 7 5 0 0 8336 0 9 4 0 0 6
709 398
709 441
938 441
938 319
917 319
917 327
5 7 6 0 0 8320 0 21 9 0 0 6
549 399
549 460
775 460
775 320
754 320
754 328
5 7 7 0 0 8320 0 14 21 0 0 6
401 395
401 403
615 403
615 321
594 321
594 329
1 6 2 0 0 4096 0 2 15 0 0 2
349 297
349 299
14 6 8 0 0 8320 0 10 5 0 0 6
657 238
657 227
805 227
805 309
820 309
820 301
14 6 9 0 0 8320 0 20 10 0 0 6
497 239
497 228
642 228
642 310
657 310
657 302
14 6 10 0 0 8320 0 15 20 0 0 6
349 235
349 225
482 225
482 311
497 311
497 303
3 1 2 0 0 4224 0 4 3 0 0 4
899 391
899 406
903 406
903 414
2 1 2 0 0 0 0 4 4 0 0 2
908 391
917 391
3 2 2 0 0 0 0 4 4 0 0 2
899 391
908 391
4 3 2 0 0 0 0 4 4 0 0 2
890 391
899 391
10 6 11 0 0 12416 0 4 4 0 0 6
863 327
863 323
849 323
849 405
863 405
863 397
2 8 12 0 0 4224 0 5 4 0 0 4
892 301
892 319
899 319
899 327
1 7 5 0 0 0 0 5 4 0 0 4
901 301
901 319
917 319
917 327
3 9 13 0 0 4224 0 5 4 0 0 4
883 301
883 319
881 319
881 327
4 10 11 0 0 0 0 5 4 0 0 4
874 301
874 319
863 319
863 327
7 7 14 0 0 8320 0 5 7 0 0 4
901 231
901 227
890 227
890 219
8 6 15 0 0 8320 0 5 7 0 0 4
892 231
892 227
884 227
884 219
9 5 16 0 0 12416 0 5 7 0 0 4
883 231
883 227
878 227
878 219
10 4 17 0 0 12416 0 5 7 0 0 4
874 231
874 227
872 227
872 219
11 3 18 0 0 12416 0 5 7 0 0 4
865 231
865 227
866 227
866 219
12 2 19 0 0 12416 0 5 7 0 0 4
856 231
856 227
860 227
860 219
13 1 20 0 0 12416 0 5 7 0 0 4
847 231
847 227
854 227
854 219
1 2 3 0 0 4224 0 6 23 0 0 2
875 88
875 99
1 9 21 0 0 4224 0 23 7 0 0 2
875 135
875 147
3 1 2 0 0 0 0 9 8 0 0 4
736 392
736 407
740 407
740 415
2 1 2 0 0 0 0 9 9 0 0 2
745 392
754 392
3 2 2 0 0 0 0 9 9 0 0 2
736 392
745 392
4 3 2 0 0 0 0 9 9 0 0 2
727 392
736 392
10 6 22 0 0 12416 0 9 9 0 0 6
700 328
700 324
686 324
686 406
700 406
700 398
2 8 23 0 0 4224 0 10 9 0 0 4
729 302
729 320
736 320
736 328
1 7 6 0 0 0 0 10 9 0 0 4
738 302
738 320
754 320
754 328
3 9 24 0 0 4224 0 10 9 0 0 4
720 302
720 320
718 320
718 328
4 10 22 0 0 0 0 10 9 0 0 4
711 302
711 320
700 320
700 328
7 7 25 0 0 8320 0 10 12 0 0 4
738 232
738 228
727 228
727 220
8 6 26 0 0 8320 0 10 12 0 0 4
729 232
729 228
721 228
721 220
9 5 27 0 0 12416 0 10 12 0 0 4
720 232
720 228
715 228
715 220
10 4 28 0 0 12416 0 10 12 0 0 4
711 232
711 228
709 228
709 220
11 3 29 0 0 12416 0 10 12 0 0 4
702 232
702 228
703 228
703 220
12 2 30 0 0 12416 0 10 12 0 0 4
693 232
693 228
697 228
697 220
13 1 31 0 0 12416 0 10 12 0 0 4
684 232
684 228
691 228
691 220
1 2 3 0 0 0 0 11 24 0 0 2
712 89
712 100
1 9 32 0 0 4224 0 24 12 0 0 2
712 136
712 148
3 1 2 0 0 0 0 14 13 0 0 4
428 389
428 404
432 404
432 412
2 1 2 0 0 0 0 14 14 0 0 2
437 389
446 389
3 2 2 0 0 0 0 14 14 0 0 2
428 389
437 389
4 3 2 0 0 0 0 14 14 0 0 2
419 389
428 389
10 6 33 0 0 12416 0 14 14 0 0 6
392 325
392 321
378 321
378 403
392 403
392 395
2 8 34 0 0 4224 0 15 14 0 0 4
421 299
421 317
428 317
428 325
1 7 35 0 0 4224 0 15 14 0 0 4
430 299
430 317
446 317
446 325
3 9 36 0 0 4224 0 15 14 0 0 4
412 299
412 317
410 317
410 325
4 10 33 0 0 0 0 15 14 0 0 4
403 299
403 317
392 317
392 325
7 7 37 0 0 8320 0 15 17 0 0 4
430 229
430 225
419 225
419 217
8 6 38 0 0 8320 0 15 17 0 0 4
421 229
421 225
413 225
413 217
9 5 39 0 0 12416 0 15 17 0 0 4
412 229
412 225
407 225
407 217
10 4 40 0 0 12416 0 15 17 0 0 4
403 229
403 225
401 225
401 217
11 3 41 0 0 12416 0 15 17 0 0 4
394 229
394 225
395 225
395 217
12 2 42 0 0 12416 0 15 17 0 0 4
385 229
385 225
389 225
389 217
13 1 43 0 0 12416 0 15 17 0 0 4
376 229
376 225
383 225
383 217
1 2 3 0 0 0 0 16 25 0 0 2
404 86
404 97
1 9 44 0 0 4224 0 25 17 0 0 2
404 133
404 145
3 1 2 0 0 0 0 21 22 0 0 4
576 393
576 408
580 408
580 416
2 1 2 0 0 0 0 21 21 0 0 2
585 393
594 393
3 2 2 0 0 0 0 21 21 0 0 2
576 393
585 393
4 3 2 0 0 0 0 21 21 0 0 2
567 393
576 393
10 6 45 0 0 12416 0 21 21 0 0 6
540 329
540 325
526 325
526 407
540 407
540 399
2 8 46 0 0 4224 0 20 21 0 0 4
569 303
569 321
576 321
576 329
1 7 7 0 0 0 0 20 21 0 0 4
578 303
578 321
594 321
594 329
3 9 47 0 0 4224 0 20 21 0 0 4
560 303
560 321
558 321
558 329
4 10 45 0 0 0 0 20 21 0 0 4
551 303
551 321
540 321
540 329
7 7 48 0 0 8320 0 20 18 0 0 4
578 233
578 229
567 229
567 221
8 6 49 0 0 8320 0 20 18 0 0 4
569 233
569 229
561 229
561 221
9 5 50 0 0 12416 0 20 18 0 0 4
560 233
560 229
555 229
555 221
10 4 51 0 0 12416 0 20 18 0 0 4
551 233
551 229
549 229
549 221
11 3 52 0 0 12416 0 20 18 0 0 4
542 233
542 229
543 229
543 221
12 2 53 0 0 12416 0 20 18 0 0 4
533 233
533 229
537 229
537 221
13 1 54 0 0 12416 0 20 18 0 0 4
524 233
524 229
531 229
531 221
1 2 3 0 0 0 0 19 26 0 0 2
552 90
552 101
1 9 55 0 0 4224 0 26 18 0 0 2
552 137
552 149
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
