CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
38 96 1497 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 96 1497 799
143654930 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 300 203 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
14 Logic Display~
6 421 387 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4441 0 0
0
0
14 Logic Display~
6 449 389 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3618 0 0
0
0
14 Logic Display~
6 475 391 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6153 0 0
0
0
14 Logic Display~
6 501 392 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5394 0 0
0
0
14 Logic Display~
6 525 392 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7734 0 0
0
0
7 Ground~
168 566 338 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9914 0 0
0
0
6 74LS83
105 651 357 0 14 29
0 13 14 15 16 10 11 12 9 2
5 6 7 8 4
0
0 0 13040 270
7 74LS83A
-24 -60 25 -52
2 U4
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3747 0 0
0
0
7 74LS273
150 371 255 0 18 37
0 3 21 10 11 12 9 17 18 19
20 13 14 15 16 10 11 12 9
0
0 0 13040 0
7 74LS273
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
3549 0 0
0
0
7 Buffer~
58 161 158 0 2 22
0 22 21
0
0 0 624 270
4 4050
-14 -19 14 -11
3 U1A
13 -5 34 3
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 1 0
1 U
7931 0 0
0
0
10 Ascii Key~
169 182 99 0 11 12
0 20 19 18 17 23 24 25 22 0
0 53
0
0 0 4656 0
0
4 KBD1
-14 -34 14 -26
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 0 0 0 0
3 KBD
9325 0 0
0
0
25
1 1 3 0 0 8320 0 1 9 0 0 4
312 203
325 203
325 219
333 219
14 1 4 0 0 8320 0 8 2 0 0 4
608 391
608 415
421 415
421 405
10 1 5 0 0 8320 0 8 3 0 0 4
662 391
662 415
449 415
449 407
11 1 6 0 0 8320 0 8 4 0 0 4
653 391
653 417
475 417
475 409
12 1 7 0 0 8320 0 8 5 0 0 4
644 391
644 418
501 418
501 410
13 1 8 0 0 8320 0 8 6 0 0 4
635 391
635 418
525 418
525 410
1 9 2 0 0 8320 0 7 8 0 0 4
566 332
566 319
608 319
608 327
18 6 9 0 0 12288 0 9 9 0 0 6
403 300
407 300
407 315
325 315
325 264
339 264
15 3 10 0 0 12288 0 9 9 0 0 6
403 273
407 273
407 199
325 199
325 237
339 237
16 4 11 0 0 8192 0 9 9 0 0 6
403 282
407 282
407 199
325 199
325 246
339 246
17 5 12 0 0 8192 0 9 9 0 0 6
403 291
407 291
407 199
325 199
325 255
339 255
11 1 13 0 0 4224 0 9 8 0 0 3
403 237
689 237
689 327
12 2 14 0 0 4224 0 9 8 0 0 3
403 246
680 246
680 327
13 3 15 0 0 4224 0 9 8 0 0 3
403 255
671 255
671 327
14 4 16 0 0 4224 0 9 8 0 0 3
403 264
662 264
662 327
15 5 10 0 0 4224 0 9 8 0 0 3
403 273
653 273
653 327
16 6 11 0 0 4224 0 9 8 0 0 3
403 282
644 282
644 327
17 7 12 0 0 4224 0 9 8 0 0 3
403 291
635 291
635 327
18 8 9 0 0 4224 0 9 8 0 0 3
403 300
626 300
626 327
4 7 17 0 0 8320 0 11 9 0 0 3
185 123
185 273
339 273
3 8 18 0 0 4224 0 11 9 0 0 3
191 123
191 282
339 282
2 9 19 0 0 4224 0 11 9 0 0 3
197 123
197 291
339 291
1 10 20 0 0 4224 0 11 9 0 0 3
203 123
203 300
339 300
2 2 21 0 0 8320 0 10 9 0 0 3
161 173
161 228
339 228
8 1 22 0 0 4224 0 11 10 0 0 2
161 123
161 143
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
