CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
38 96 1497 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 96 1497 799
143654930 0
0
6 Title:
5 Name:
0
0
0
22
14 Logic Display~
6 611 419 0 1 2
10 0
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L3
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8953 0 0
0
0
14 Logic Display~
6 632 419 0 1 2
10 0
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L2
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4441 0 0
0
0
14 Logic Display~
6 650 421 0 1 2
10 0
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L1
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3618 0 0
0
0
7 Pulser~
4 159 311 0 8 12
0 0 0 0 0 0 0 5 5
0
0 0 4640 0
0
2 V6
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 326 472 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 175 423 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
7734 0 0
0
0
9 2-In AND~
219 323 355 0 1 22
0 0
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 2065446846
65 0 0 0 4 1 3 0
1 U
9914 0 0
0
0
8 2-In OR~
219 423 368 0 1 22
0 0
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U6A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 1746679725
65 0 0 0 4 1 2 0
1 U
3747 0 0
0
0
13 Logic Switch~
5 416 256 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3549 0 0
0
0
7 Ground~
168 676 315 0 1 3
0 0
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7931 0 0
0
0
6 74LS93
109 560 347 0 1 17
0 0
0
0 0 13024 0
6 74LS93
-21 -35 21 -27
2 U5
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
9325 0 0
0
0
7 Ground~
168 789 252 0 1 3
0 0
0
0 0 53344 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8903 0 0
0
0
13 Logic Switch~
5 1141 483 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 21344 512
2 5V
-7 -16 7 -8
2 V1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3834 0 0
0
0
6 1K RAM
79 736 322 0 1 41
0 0
0
0 0 13024 0
5 RAM1K
-17 -19 18 -11
2 U4
-7 -70 7 -62
0
15 DVCC=22;DGND=11
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 0 0 0 0 0
1 U
3363 0 0
0
0
7 Ground~
168 1175 266 0 1 3
0 0
0
0 0 53344 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7668 0 0
0
0
7 Buffer~
58 1234 318 0 2 22
0 30 29
0
0 0 608 180
4 4050
-14 -19 14 -11
3 U1A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 1 0
1 U
4718 0 0
0
0
10 Ascii Key~
169 1298 342 0 11 12
0 28 27 26 25 40 41 42 30 0
0 56
0
0 0 4640 270
0
4 KBD1
-12 -38 16 -30
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
3874 0 0
0
0
7 74LS173
129 1116 323 0 1 29
0 0
0
0 0 13024 512
7 74LS173
-24 -51 25 -43
2 U3
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
6671 0 0
0
0
9 Resistor~
219 922 97 0 4 5
0 38 3 0 1
0
0 0 864 90
3 330
5 0 26 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3789 0 0
0
0
6 74LS47
187 907 244 0 14 29
0 15 14 13 12 44 45 31 32 33
34 35 36 37 46
0
0 0 13024 602
6 74LS47
-21 -60 21 -52
2 U2
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
4871 0 0
0
0
2 +V
167 922 59 0 1 3
0 3
0
0 0 54240 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3750 0 0
0
0
9 CA 7-Seg~
184 922 163 0 18 19
10 37 36 35 34 33 32 31 43 38
0 2 0 0 2 0 0 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
8778 0 0
0
0
50
1 0 0 0 0 0 0 1 0 0 18 4
611 405
611 343
612 343
612 338
1 0 0 0 0 0 0 2 0 0 19 2
632 405
632 347
1 0 0 0 0 0 0 3 0 0 20 4
650 407
650 361
651 361
651 356
3 1 0 0 0 0 0 4 7 0 0 4
183 302
291 302
291 346
299 346
1 2 0 0 0 0 0 6 7 0 0 4
187 423
291 423
291 364
299 364
3 1 0 0 0 0 0 7 8 0 0 4
344 355
402 355
402 359
410 359
1 2 0 0 0 0 0 5 8 0 0 4
338 472
402 472
402 377
410 377
3 4 0 0 0 0 0 8 11 0 0 4
456 368
514 368
514 365
522 365
1 2 0 0 0 0 0 9 11 0 0 4
428 256
514 256
514 347
528 347
1 1 0 0 0 0 0 9 11 0 0 4
428 256
514 256
514 338
528 338
1 0 0 0 0 0 0 10 0 0 16 4
676 309
676 301
696 301
696 296
6 0 0 0 0 0 0 14 0 0 17 3
704 331
704 332
696 332
5 0 0 0 0 0 0 14 0 0 17 3
704 322
704 320
696 320
4 0 0 0 0 0 0 14 0 0 17 3
704 313
704 314
696 314
3 0 0 0 0 0 0 14 0 0 17 3
704 304
704 305
696 305
2 0 0 0 0 0 0 14 0 0 17 3
704 295
704 296
696 296
7 1 0 0 0 0 0 14 14 0 0 4
704 340
696 340
696 286
704 286
5 8 0 0 0 0 0 11 14 0 0 4
592 338
696 338
696 349
704 349
6 9 0 0 0 0 0 11 14 0 0 4
592 347
696 347
696 358
704 358
7 10 0 0 0 0 0 11 14 0 0 4
592 356
696 356
696 367
704 367
19 1 0 0 0 0 0 14 12 0 0 3
774 286
789 286
789 260
1 0 0 0 0 0 0 20 0 0 26 2
948 281
948 340
2 0 0 0 0 0 0 20 0 0 27 2
939 281
939 349
3 0 0 0 0 0 0 20 0 0 28 2
930 281
930 358
4 0 0 0 0 0 0 20 0 0 29 4
921 281
921 362
922 362
922 367
15 11 0 0 0 0 0 14 18 0 0 4
768 340
1070 340
1070 332
1084 332
16 12 0 0 0 0 0 14 18 0 0 4
768 349
1070 349
1070 341
1084 341
17 13 0 0 0 0 0 14 18 0 0 4
768 358
1070 358
1070 350
1084 350
18 14 0 0 0 0 0 14 18 0 0 4
768 367
1070 367
1070 359
1084 359
10 0 0 0 0 0 0 18 0 0 32 3
1078 305
1078 307
991 307
9 0 0 0 0 0 0 18 0 0 32 3
1078 296
1078 295
991 295
20 1 0 0 0 0 0 14 13 0 0 4
774 295
991 295
991 483
1129 483
3 0 0 0 0 0 0 18 0 0 34 3
1154 314
1175 314
1175 277
2 0 0 0 0 0 0 18 0 0 35 4
1154 305
1170 305
1170 277
1175 277
1 1 0 0 0 0 0 18 15 0 0 3
1148 296
1175 296
1175 274
5 4 0 0 0 0 0 18 17 0 0 4
1148 332
1266 332
1266 345
1274 345
6 3 0 0 0 0 0 18 17 0 0 4
1148 341
1266 341
1266 351
1274 351
7 2 0 0 0 0 0 18 17 0 0 4
1148 350
1266 350
1266 357
1274 357
8 1 0 0 0 0 0 18 17 0 0 4
1148 359
1266 359
1266 363
1274 363
4 2 0 0 0 0 0 18 16 0 0 4
1148 323
1211 323
1211 318
1219 318
1 8 0 0 0 0 0 16 17 0 0 4
1249 318
1266 318
1266 321
1274 321
7 7 31 0 0 0 0 20 22 0 0 4
948 211
948 207
937 207
937 199
8 6 32 0 0 0 0 20 22 0 0 4
939 211
939 207
931 207
931 199
9 5 33 0 0 0 0 20 22 0 0 4
930 211
930 207
925 207
925 199
10 4 34 0 0 0 0 20 22 0 0 4
921 211
921 207
919 207
919 199
11 3 35 0 0 0 0 20 22 0 0 4
912 211
912 207
913 207
913 199
12 2 36 0 0 0 0 20 22 0 0 4
903 211
903 207
907 207
907 199
13 1 37 0 0 0 0 20 22 0 0 4
894 211
894 207
901 207
901 199
1 2 3 0 0 0 0 21 19 0 0 2
922 68
922 79
1 9 38 0 0 0 0 19 22 0 0 2
922 115
922 127
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
301 477 333 501
311 485 335 501
3 SW3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
150 433 182 457
160 441 184 457
3 SW2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
338 240 370 264
348 248 372 264
3 SW1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1157 461 1189 485
1167 469 1191 485
3 SW4
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
