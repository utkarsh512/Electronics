CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 2 100 9
38 96 1497 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 96 1497 799
143654930 0
0
6 Title:
5 Name:
0
0
0
29
13 Logic Switch~
5 326 472 0 1 11
0 28
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 175 423 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 416 256 0 1 11
0 30
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 1141 483 0 10 11
0 31 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6153 0 0
0
0
7 Ground~
168 374 164 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5394 0 0
0
0
7 74LS138
19 339 97 0 14 29
0 13 12 11 38 2 2 14 15 16
17 18 19 20 21
0
0 0 13296 90
7 74LS138
52 -3 101 5
2 U8
70 -13 84 -5
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 512 1 0 0 0
1 U
7734 0 0
0
0
6 74LS48
188 910 237 0 14 29
0 22 23 24 25 39 3 4 5 6
7 8 9 10 3
0
0 0 13040 602
6 74LS48
-21 -60 21 -52
2 U2
57 -3 71 5
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
9914 0 0
0
0
9 CC 7-Seg~
183 1184 103 0 18 19
10 10 9 8 7 6 5 4 40 14
0 0 0 0 0 0 0 2 1
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP8
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3747 0 0
0
0
9 CC 7-Seg~
183 1081 103 0 18 19
10 10 9 8 7 6 5 4 41 15
0 0 0 0 0 0 0 2 1
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP7
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3549 0 0
0
0
9 CC 7-Seg~
183 974 103 0 17 19
10 10 9 8 7 6 5 4 42 16
0 0 0 0 0 0 0 2
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP6
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
7931 0 0
0
0
9 CC 7-Seg~
183 873 102 0 18 19
10 10 9 8 7 6 5 4 43 17
0 0 0 0 0 0 0 2 1
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP5
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
9325 0 0
0
0
9 CC 7-Seg~
183 774 103 0 18 19
10 10 9 8 7 6 5 4 44 18
0 0 0 0 0 0 0 2 1
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP4
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
8903 0 0
0
0
9 CC 7-Seg~
183 675 103 0 18 19
10 10 9 8 7 6 5 4 45 19
0 0 0 0 0 0 0 2 1
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP3
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3834 0 0
0
0
9 CC 7-Seg~
183 576 104 0 18 19
10 10 9 8 7 6 5 4 46 20
0 0 0 0 0 0 0 2 1
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3363 0 0
0
0
9 CC 7-Seg~
183 470 105 0 18 19
10 10 9 8 7 6 5 4 47 21
0 0 0 0 0 0 0 2 1
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
7668 0 0
0
0
14 Logic Display~
6 611 419 0 1 2
10 13
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L3
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4718 0 0
0
0
14 Logic Display~
6 632 419 0 1 2
10 12
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L2
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3874 0 0
0
0
14 Logic Display~
6 650 421 0 1 2
10 11
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L1
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6671 0 0
0
0
7 Pulser~
4 159 311 0 10 12
0 48 49 3 50 0 0 5 5 2
7
0
0 0 4656 0
0
2 V6
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3789 0 0
0
0
9 2-In AND~
219 323 355 0 3 22
0 3 26 27
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 2065446846
65 0 0 0 4 1 3 0
1 U
4871 0 0
0
0
8 2-In OR~
219 423 368 0 3 22
0 27 28 29
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U6A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 1746679725
65 0 0 0 4 1 2 0
1 U
3750 0 0
0
0
7 Ground~
168 676 315 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8778 0 0
0
0
6 74LS93
109 560 347 0 8 17
0 30 30 51 29 13 12 11 52
0
0 0 13040 0
6 74LS93
-21 -35 21 -27
2 U5
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 512 1 0 0 0
1 U
538 0 0
0
0
7 Ground~
168 789 252 0 1 3
0 2
0
0 0 53360 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6843 0 0
0
0
6 1K RAM
79 736 322 0 20 41
0 2 2 2 2 2 2 2 13 12
11 53 54 55 56 22 23 24 25 2
31
0
0 0 13040 0
5 RAM1K
-17 -19 18 -11
2 U4
-7 -70 7 -62
0
15 DVCC=22;DGND=11
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 512 1 0 0 0
1 U
3136 0 0
0
0
7 Ground~
168 1175 266 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5950 0 0
0
0
7 Buffer~
58 1234 318 0 2 22
0 37 36
0
0 0 624 180
4 4050
-14 -19 14 -11
3 U1A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 1 0
1 U
5670 0 0
0
0
10 Ascii Key~
169 1298 342 0 11 12
0 35 34 33 32 57 58 59 37 0
0 56
0
0 0 4656 270
0
4 KBD1
-12 -38 16 -30
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
6828 0 0
0
0
7 74LS173
129 1116 323 0 14 29
0 2 2 2 36 32 33 34 35 31
31 22 23 24 25
0
0 0 13040 512
7 74LS173
-24 -51 25 -43
2 U3
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
6735 0 0
0
0
112
0 6 3 0 0 4096 0 0 7 2 0 4
837 199
837 279
867 279
867 271
3 14 3 0 0 4224 0 19 7 0 0 5
183 302
700 302
700 199
867 199
867 207
7 7 4 0 0 4096 0 7 8 0 0 3
948 207
1199 207
1199 139
7 7 4 0 0 0 0 7 9 0 0 4
948 207
948 202
1096 202
1096 139
7 7 4 0 0 0 0 7 10 0 0 4
948 207
948 195
989 195
989 139
7 7 4 0 0 0 0 7 11 0 0 4
948 207
948 184
888 184
888 138
7 7 4 0 0 0 0 7 12 0 0 4
948 207
948 178
789 178
789 139
7 7 4 0 0 8192 0 7 13 0 0 4
948 207
948 171
690 171
690 139
7 7 4 0 0 8192 0 7 14 0 0 4
948 207
948 164
591 164
591 140
7 7 4 0 0 8320 0 7 15 0 0 4
948 207
948 157
485 157
485 141
8 6 5 0 0 8192 0 7 8 0 0 4
939 207
939 188
1193 188
1193 139
8 6 5 0 0 16 0 7 9 0 0 4
939 207
939 180
1090 180
1090 139
8 6 5 0 0 0 0 7 10 0 0 4
939 207
939 147
983 147
983 139
8 6 5 0 0 0 0 7 11 0 0 4
939 207
939 146
882 146
882 138
8 6 5 0 0 0 0 7 12 0 0 4
939 207
939 147
783 147
783 139
8 6 5 0 0 8192 0 7 13 0 0 4
939 207
939 147
684 147
684 139
8 6 5 0 0 8192 0 7 14 0 0 4
939 207
939 148
585 148
585 140
8 6 5 0 0 8320 0 7 15 0 0 4
939 207
939 149
479 149
479 141
9 5 6 0 0 8192 0 7 8 0 0 4
930 207
930 147
1187 147
1187 139
9 5 6 0 0 0 0 7 9 0 0 4
930 207
930 147
1084 147
1084 139
9 5 6 0 0 0 0 7 10 0 0 4
930 207
930 147
977 147
977 139
9 5 6 0 0 0 0 7 11 0 0 4
930 207
930 146
876 146
876 138
9 5 6 0 0 0 0 7 12 0 0 4
930 207
930 147
777 147
777 139
9 5 6 0 0 0 0 7 13 0 0 4
930 207
930 147
678 147
678 139
9 5 6 0 0 8192 0 7 14 0 0 4
930 207
930 148
579 148
579 140
9 5 6 0 0 8320 0 7 15 0 0 4
930 207
930 149
473 149
473 141
10 4 7 0 0 8192 0 7 8 0 0 4
921 207
921 147
1181 147
1181 139
10 4 7 0 0 0 0 7 9 0 0 4
921 207
921 147
1078 147
1078 139
10 4 7 0 0 0 0 7 10 0 0 4
921 207
921 147
971 147
971 139
10 4 7 0 0 0 0 7 11 0 0 4
921 207
921 146
870 146
870 138
10 4 7 0 0 0 0 7 12 0 0 4
921 207
921 147
771 147
771 139
10 4 7 0 0 0 0 7 13 0 0 4
921 207
921 147
672 147
672 139
10 4 7 0 0 8192 0 7 14 0 0 4
921 207
921 148
573 148
573 140
10 4 7 0 0 8320 0 7 15 0 0 4
921 207
921 149
467 149
467 141
11 3 8 0 0 8192 0 7 8 0 0 4
912 207
912 147
1175 147
1175 139
11 3 8 0 0 0 0 7 9 0 0 4
912 207
912 147
1072 147
1072 139
11 3 8 0 0 0 0 7 10 0 0 4
912 207
912 147
965 147
965 139
11 3 8 0 0 0 0 7 11 0 0 4
912 207
912 146
864 146
864 138
11 3 8 0 0 0 0 7 12 0 0 4
912 207
912 147
765 147
765 139
11 3 8 0 0 0 0 7 13 0 0 4
912 207
912 147
666 147
666 139
11 3 8 0 0 8192 0 7 14 0 0 4
912 207
912 148
567 148
567 140
11 3 8 0 0 8320 0 7 15 0 0 4
912 207
912 149
461 149
461 141
12 2 9 0 0 8192 0 7 8 0 0 4
903 207
903 147
1169 147
1169 139
12 2 9 0 0 0 0 7 9 0 0 4
903 207
903 147
1066 147
1066 139
12 2 9 0 0 0 0 7 10 0 0 4
903 207
903 147
959 147
959 139
12 2 9 0 0 0 0 7 11 0 0 4
903 207
903 146
858 146
858 138
12 2 9 0 0 0 0 7 12 0 0 4
903 207
903 147
759 147
759 139
12 2 9 0 0 0 0 7 13 0 0 4
903 207
903 147
660 147
660 139
12 2 9 0 0 8192 0 7 14 0 0 4
903 207
903 148
561 148
561 140
12 2 9 0 0 8320 0 7 15 0 0 4
903 207
903 149
455 149
455 141
13 1 10 0 0 8192 0 7 8 0 0 4
894 207
894 147
1163 147
1163 139
13 1 10 0 0 0 0 7 9 0 0 4
894 207
894 147
1060 147
1060 139
13 1 10 0 0 0 0 7 10 0 0 4
894 207
894 147
953 147
953 139
13 1 10 0 0 0 0 7 11 0 0 4
894 207
894 146
852 146
852 138
13 1 10 0 0 0 0 7 12 0 0 4
894 207
894 147
753 147
753 139
13 1 10 0 0 0 0 7 13 0 0 4
894 207
894 147
654 147
654 139
13 1 10 0 0 8192 0 7 14 0 0 4
894 207
894 148
555 148
555 140
13 1 10 0 0 8320 0 7 15 0 0 4
894 207
894 149
449 149
449 141
6 1 2 0 0 4096 0 6 5 0 0 4
378 132
378 150
374 150
374 158
5 1 2 0 0 0 0 6 5 0 0 4
369 132
369 150
374 150
374 158
3 0 11 0 0 8320 0 6 0 0 95 4
333 126
333 277
654 277
654 356
2 0 12 0 0 8320 0 6 0 0 77 5
324 126
324 291
627 291
627 349
632 349
1 0 13 0 0 8320 0 6 0 0 76 5
315 126
315 316
607 316
607 338
612 338
7 9 14 0 0 8320 0 6 8 0 0 4
315 56
315 5
1184 5
1184 61
8 9 15 0 0 8320 0 6 9 0 0 4
324 56
324 10
1081 10
1081 61
9 9 16 0 0 8320 0 6 10 0 0 4
333 56
333 15
974 15
974 61
10 9 17 0 0 8320 0 6 11 0 0 4
342 56
342 19
873 19
873 60
11 9 18 0 0 8320 0 6 12 0 0 4
351 56
351 24
774 24
774 61
12 9 19 0 0 8320 0 6 13 0 0 4
360 56
360 30
675 30
675 61
13 9 20 0 0 8320 0 6 14 0 0 4
369 56
369 37
576 37
576 62
14 9 21 0 0 8320 0 6 15 0 0 4
378 56
378 45
470 45
470 63
1 0 22 0 0 4096 0 7 0 0 97 2
948 271
948 340
2 0 23 0 0 4096 0 7 0 0 98 4
939 271
939 344
940 344
940 349
3 0 24 0 0 4096 0 7 0 0 99 2
930 271
930 358
4 0 25 0 0 4096 0 7 0 0 100 4
921 271
921 362
922 362
922 367
1 0 13 0 0 0 0 16 0 0 93 4
611 405
611 343
612 343
612 338
1 0 12 0 0 0 0 17 0 0 94 2
632 405
632 347
1 0 11 0 0 0 0 18 0 0 95 4
650 407
650 361
651 361
651 356
3 1 3 0 0 128 0 19 20 0 0 4
183 302
291 302
291 346
299 346
1 2 26 0 0 4224 0 2 20 0 0 4
187 423
291 423
291 364
299 364
3 1 27 0 0 4224 0 20 21 0 0 4
344 355
402 355
402 359
410 359
1 2 28 0 0 8320 0 1 21 0 0 4
338 472
402 472
402 377
410 377
3 4 29 0 0 4224 0 21 23 0 0 4
456 368
514 368
514 365
522 365
1 2 30 0 0 8320 0 3 23 0 0 4
428 256
514 256
514 347
528 347
1 1 30 0 0 0 0 3 23 0 0 4
428 256
514 256
514 338
528 338
1 0 2 0 0 8192 0 22 0 0 91 4
676 309
676 301
696 301
696 296
6 0 2 0 0 0 0 25 0 0 92 3
704 331
704 332
696 332
5 0 2 0 0 0 0 25 0 0 92 3
704 322
704 320
696 320
4 0 2 0 0 0 0 25 0 0 92 3
704 313
704 314
696 314
3 0 2 0 0 0 0 25 0 0 92 3
704 304
704 305
696 305
2 0 2 0 0 0 0 25 0 0 92 3
704 295
704 296
696 296
7 1 2 0 0 8320 0 25 25 0 0 4
704 340
696 340
696 286
704 286
5 8 13 0 0 128 0 23 25 0 0 4
592 338
696 338
696 349
704 349
6 9 12 0 0 128 0 23 25 0 0 4
592 347
696 347
696 358
704 358
7 10 11 0 0 128 0 23 25 0 0 4
592 356
696 356
696 367
704 367
19 1 2 0 0 0 0 25 24 0 0 3
774 286
789 286
789 260
15 11 22 0 0 4224 0 25 29 0 0 4
768 340
1070 340
1070 332
1084 332
16 12 23 0 0 4224 0 25 29 0 0 4
768 349
1070 349
1070 341
1084 341
17 13 24 0 0 4224 0 25 29 0 0 4
768 358
1070 358
1070 350
1084 350
18 14 25 0 0 4224 0 25 29 0 0 4
768 367
1070 367
1070 359
1084 359
10 0 31 0 0 8192 0 29 0 0 103 3
1078 305
1078 307
991 307
9 0 31 0 0 0 0 29 0 0 103 3
1078 296
1078 295
991 295
20 1 31 0 0 4224 0 25 4 0 0 4
774 295
991 295
991 483
1129 483
3 0 2 0 0 0 0 29 0 0 105 3
1154 314
1175 314
1175 277
2 0 2 0 0 0 0 29 0 0 106 4
1154 305
1170 305
1170 277
1175 277
1 1 2 0 0 0 0 29 26 0 0 3
1148 296
1175 296
1175 274
5 4 32 0 0 4224 0 29 28 0 0 4
1148 332
1266 332
1266 345
1274 345
6 3 33 0 0 4224 0 29 28 0 0 4
1148 341
1266 341
1266 351
1274 351
7 2 34 0 0 4224 0 29 28 0 0 4
1148 350
1266 350
1266 357
1274 357
8 1 35 0 0 4224 0 29 28 0 0 4
1148 359
1266 359
1266 363
1274 363
4 2 36 0 0 4224 0 29 27 0 0 4
1148 323
1211 323
1211 318
1219 318
1 8 37 0 0 4224 0 27 28 0 0 4
1249 318
1266 318
1266 321
1274 321
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
444 180 524 204
454 188 526 204
9 18EC30048
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1157 461 1189 485
1167 469 1191 485
3 SW4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
338 240 370 264
348 248 372 264
3 SW1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
150 433 182 457
160 441 184 457
3 SW2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
301 477 333 501
311 485 335 501
3 SW3
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
