CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
20 0 23 130 9
38 96 1497 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 96 1497 799
143654930 0
0
6 Title:
5 Name:
0
0
0
29
13 Logic Switch~
5 75 238 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 610 98 0 1 11
0 8
0
0 0 21360 512
2 0V
-7 -16 7 -8
2 V5
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 394 255 0 1 11
0 7
0
0 0 21360 512
2 0V
-7 -16 7 -8
2 V4
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 401 19 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
9 2-In AND~
219 483 296 0 3 22
0 6 5 4
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 299108277
65 0 0 0 4 2 1 0
1 U
5394 0 0
0
0
9 Inverter~
13 400 295 0 2 22
0 7 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U11C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 3 3 0
1 U
7734 0 0
0
0
9 Inverter~
13 335 145 0 2 22
0 15 14
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U11B
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 3 0
1 U
9914 0 0
0
0
7 Ground~
168 310 329 0 1 3
0 2
0
0 0 53360 180
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3747 0 0
0
0
8 2-In OR~
219 382 182 0 3 22
0 14 5 29
0
0 0 624 782
6 74LS32
-21 -24 21 -16
4 U10A
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 349505457
65 0 0 0 4 1 2 0
1 U
3549 0 0
0
0
9 2-In AND~
219 352 247 0 3 22
0 7 29 28
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U9A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 366282672
65 0 0 0 4 1 1 0
1 U
7931 0 0
0
0
7 Ground~
168 342 338 0 1 3
0 2
0
0 0 53360 180
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9325 0 0
0
0
7 Ground~
168 176 92 0 1 3
0 2
0
0 0 53360 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8903 0 0
0
0
7 Ground~
168 42 93 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3834 0 0
0
0
8 Hex Key~
166 232 61 0 11 12
0 43 44 45 46 0 0 0 0 0
15 70
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3363 0 0
0
0
8 Hex Key~
166 86 62 0 11 12
0 47 48 49 50 0 0 0 0 0
2 50
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
7668 0 0
0
0
6 74LS93
109 632 177 0 8 17
0 8 8 4 19 16 17 18 19
0
0 0 13040 782
6 74LS93
-21 -35 21 -27
2 U8
28 0 42 8
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
4718 0 0
0
0
6 74LS83
105 300 390 0 14 29
0 9 10 11 12 2 67 68 2 2
23 22 21 20 30
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
2 U7
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3874 0 0
0
0
6 74LS83
105 151 390 0 14 29
0 34 33 32 31 69 70 71 72 30
27 26 25 24 5
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
2 U6
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
6671 0 0
0
0
7 74LS273
150 167 268 0 18 37
0 13 28 42 41 40 39 38 37 36
35 34 33 32 31 9 10 11 12
0
0 0 13040 782
7 74LS273
-24 -60 25 -52
2 U5
54 0 68 8
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
3789 0 0
0
0
7 74LS157
122 93 154 0 14 29
0 15 24 47 25 48 26 49 27 50
2 39 40 41 42
0
0 0 13040 270
7 74LS157
-24 -60 25 -52
2 U2
54 0 68 8
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
4871 0 0
0
0
7 74LS157
122 232 153 0 14 29
0 15 20 43 21 44 22 45 23 46
2 35 36 37 38
0
0 0 13040 270
7 74LS157
-24 -60 25 -52
2 U3
54 0 68 8
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3750 0 0
0
0
6 74LS47
187 1016 223 0 14 29
0 9 10 11 12 73 74 59 60 61
62 63 64 65 75
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U4
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
8778 0 0
0
0
2 +V
167 1031 38 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
538 0 0
0
0
9 CA 7-Seg~
184 1031 142 0 18 19
10 65 64 63 62 61 60 59 76 66
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
6843 0 0
0
0
9 CA 7-Seg~
184 883 138 0 18 19
10 57 56 55 54 53 52 51 77 58
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3136 0 0
0
0
2 +V
167 883 34 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5950 0 0
0
0
6 74LS47
187 868 219 0 14 29
0 16 17 18 19 78 79 51 52 53
54 55 56 57 80
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U1
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
5670 0 0
0
0
9 Resistor~
219 1031 76 0 4 5
0 66 3 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6828 0 0
0
0
9 Resistor~
219 883 72 0 4 5
0 58 3 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6735 0 0
0
0
80
3 3 4 0 0 8320 0 5 16 0 0 5
504 296
661 296
661 135
637 135
637 143
14 2 5 0 0 8192 0 18 5 0 0 5
194 424
194 428
451 428
451 305
459 305
2 1 6 0 0 4224 0 6 5 0 0 4
421 295
451 295
451 287
459 287
1 1 7 0 0 8320 0 3 6 0 0 4
382 255
377 255
377 295
385 295
1 0 8 0 0 8320 0 2 0 0 6 5
598 98
596 98
596 144
622 144
622 149
1 2 8 0 0 0 0 16 16 0 0 2
619 149
628 149
15 1 9 0 0 8320 0 19 22 0 0 4
180 305
180 311
1057 311
1057 260
16 2 10 0 0 8320 0 19 22 0 0 4
189 305
189 311
1048 311
1048 260
17 3 11 0 0 8320 0 19 22 0 0 4
198 305
198 311
1039 311
1039 260
18 4 12 0 0 8320 0 19 22 0 0 4
207 305
207 311
1030 311
1030 260
1 1 13 0 0 4224 0 1 19 0 0 5
87 238
107 238
107 233
126 233
126 235
2 1 14 0 0 8320 0 7 9 0 0 4
338 163
338 161
376 161
376 166
1 1 15 0 0 8192 0 4 7 0 0 3
389 19
338 19
338 127
5 1 16 0 0 8320 0 16 27 0 0 4
619 213
619 264
909 264
909 256
6 2 17 0 0 8320 0 16 27 0 0 4
628 213
628 264
900 264
900 256
7 3 18 0 0 8320 0 16 27 0 0 4
637 213
637 264
891 264
891 256
8 4 19 0 0 8320 0 16 27 0 0 4
646 213
646 264
882 264
882 256
13 2 20 0 0 12416 0 17 21 0 0 6
316 424
316 462
556 462
556 107
258 107
258 126
4 12 21 0 0 12416 0 21 17 0 0 6
240 126
240 102
563 102
563 466
307 466
307 424
6 11 22 0 0 12416 0 21 17 0 0 6
222 126
222 99
568 99
568 471
298 471
298 424
10 8 23 0 0 12416 0 17 21 0 0 6
289 424
289 475
574 475
574 95
204 95
204 126
13 2 24 0 0 12416 0 18 20 0 0 6
167 424
167 438
10 438
10 105
119 105
119 127
12 4 25 0 0 12416 0 18 20 0 0 6
158 424
158 433
17 433
17 109
101 109
101 127
11 6 26 0 0 12416 0 18 20 0 0 6
149 424
149 428
22 428
22 113
83 113
83 127
10 8 27 0 0 12416 0 18 20 0 0 6
140 424
140 423
29 423
29 117
65 117
65 127
8 0 2 0 0 4224 0 17 0 0 27 3
325 360
325 341
310 341
5 1 2 0 0 0 0 17 8 0 0 4
298 360
298 345
310 345
310 337
8 4 19 0 0 0 0 16 16 0 0 6
646 213
646 210
730 210
730 128
646 128
646 143
2 3 28 0 0 8320 0 19 10 0 0 5
135 241
135 231
319 231
319 247
325 247
1 1 7 0 0 0 0 3 10 0 0 4
382 255
380 255
380 256
370 256
3 2 29 0 0 4224 0 9 10 0 0 3
385 212
385 238
370 238
14 2 5 0 0 8320 0 18 9 0 0 6
194 424
194 443
549 443
549 147
394 147
394 166
1 9 2 0 0 0 0 11 17 0 0 4
342 346
342 352
343 352
343 360
14 9 30 0 0 8320 0 17 18 0 0 6
343 424
343 436
223 436
223 359
194 359
194 360
1 1 15 0 0 8192 0 21 4 0 0 4
267 126
267 114
389 114
389 19
1 1 15 0 0 8320 0 20 4 0 0 5
128 127
128 14
387 14
387 19
389 19
1 10 2 0 0 0 0 12 21 0 0 4
176 100
176 112
186 112
186 120
1 10 2 0 0 0 0 13 20 0 0 4
42 101
42 113
47 113
47 121
18 4 12 0 0 0 0 19 17 0 0 4
207 305
207 315
289 315
289 360
17 3 11 0 0 0 0 19 17 0 0 4
198 305
198 325
280 325
280 360
16 2 10 0 0 0 0 19 17 0 0 4
189 305
189 341
271 341
271 360
15 1 9 0 0 0 0 19 17 0 0 4
180 305
180 352
262 352
262 360
14 4 31 0 0 4224 0 19 18 0 0 4
171 305
171 352
140 352
140 360
13 3 32 0 0 4224 0 19 18 0 0 4
162 305
162 340
131 340
131 360
12 2 33 0 0 8320 0 19 18 0 0 4
153 305
153 329
122 329
122 360
11 1 34 0 0 12416 0 19 18 0 0 4
144 305
144 319
113 319
113 360
11 10 35 0 0 8320 0 21 19 0 0 4
249 190
249 227
207 227
207 241
12 9 36 0 0 8320 0 21 19 0 0 4
231 190
231 215
198 215
198 241
13 8 37 0 0 12416 0 21 19 0 0 4
213 190
213 211
189 211
189 241
14 7 38 0 0 12416 0 21 19 0 0 4
195 190
195 203
180 203
180 241
11 6 39 0 0 8320 0 20 19 0 0 4
110 191
110 201
171 201
171 241
12 5 40 0 0 8320 0 20 19 0 0 4
92 191
92 208
162 208
162 241
13 4 41 0 0 8320 0 20 19 0 0 4
74 191
74 217
153 217
153 241
14 3 42 0 0 8320 0 20 19 0 0 4
56 191
56 227
144 227
144 241
1 3 43 0 0 4224 0 14 21 0 0 4
241 85
241 112
249 112
249 126
2 5 44 0 0 4224 0 14 21 0 0 4
235 85
235 112
231 112
231 126
3 7 45 0 0 12416 0 14 21 0 0 4
229 85
229 98
213 98
213 126
4 9 46 0 0 12416 0 14 21 0 0 4
223 85
223 94
195 94
195 126
1 3 47 0 0 12416 0 15 20 0 0 4
95 86
95 99
110 99
110 127
2 5 48 0 0 12416 0 15 20 0 0 4
89 86
89 105
92 105
92 127
3 7 49 0 0 12416 0 15 20 0 0 4
83 86
83 105
74 105
74 127
4 9 50 0 0 12416 0 15 20 0 0 4
77 86
77 97
56 97
56 127
7 7 51 0 0 8320 0 27 25 0 0 4
909 186
909 182
898 182
898 174
8 6 52 0 0 8320 0 27 25 0 0 4
900 186
900 182
892 182
892 174
9 5 53 0 0 12416 0 27 25 0 0 4
891 186
891 182
886 182
886 174
10 4 54 0 0 12416 0 27 25 0 0 4
882 186
882 182
880 182
880 174
11 3 55 0 0 12416 0 27 25 0 0 4
873 186
873 182
874 182
874 174
12 2 56 0 0 12416 0 27 25 0 0 4
864 186
864 182
868 182
868 174
13 1 57 0 0 12416 0 27 25 0 0 4
855 186
855 182
862 182
862 174
1 2 3 0 0 4224 0 26 29 0 0 2
883 43
883 54
1 9 58 0 0 4224 0 29 25 0 0 2
883 90
883 102
7 7 59 0 0 8320 0 22 24 0 0 4
1057 190
1057 186
1046 186
1046 178
8 6 60 0 0 8320 0 22 24 0 0 4
1048 190
1048 186
1040 186
1040 178
9 5 61 0 0 12416 0 22 24 0 0 4
1039 190
1039 186
1034 186
1034 178
10 4 62 0 0 12416 0 22 24 0 0 4
1030 190
1030 186
1028 186
1028 178
11 3 63 0 0 12416 0 22 24 0 0 4
1021 190
1021 186
1022 186
1022 178
12 2 64 0 0 12416 0 22 24 0 0 4
1012 190
1012 186
1016 186
1016 178
13 1 65 0 0 12416 0 22 24 0 0 4
1003 190
1003 186
1010 186
1010 178
1 2 3 0 0 0 0 23 28 0 0 2
1031 47
1031 58
1 9 66 0 0 4224 0 28 24 0 0 2
1031 94
1031 106
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
408 8 464 32
415 14 463 30
6 select
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
624 81 672 105
632 87 672 103
5 reset
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
401 242 433 266
409 248 433 264
3 clk
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
