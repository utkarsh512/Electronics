CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
38 96 1497 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 96 1497 799
143654930 0
0
6 Title:
5 Name:
0
0
0
16
13 Logic Switch~
5 300 203 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
11 2-Input OR~
1 689 619 0 3 22
0 5 6 4
0
0 0 880 0
6 74LS32
-13 -25 29 -17
3 U5B
-3 -35 18 -27
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 -151380536
65 0 0 0 4 2 2 0
1 U
4441 0 0
0
0
12 2-Input AND~
0 667 557 0 3 22
0 8 7 5
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U6A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -419750439
65 0 0 0 4 1 3 0
1 U
3618 0 0
0
0
11 2-Input OR~
1 647 477 0 3 22
0 9 10 7
0
0 0 880 270
6 74LS32
29 -2 71 6
3 U5A
39 -12 60 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -151380536
65 0 0 0 4 1 2 0
1 U
6153 0 0
0
0
7 Ground~
168 832 501 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5394 0 0
0
0
14 Logic Display~
6 945 130 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7734 0 0
0
0
6 74LS83
105 875 436 0 14 29
0 8 9 10 11 2 4 4 2 2
15 14 13 12 44
0
0 0 13040 0
7 74LS83A
-24 -60 25 -52
2 U7
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
9914 0 0
0
0
7 Ground~
168 566 338 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3747 0 0
0
0
6 74LS83
105 651 357 0 14 29
0 21 22 23 24 18 19 20 17 2
8 9 10 11 6
0
0 0 13040 270
7 74LS83A
-24 -60 25 -52
2 U4
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3549 0 0
0
0
7 74LS273
150 371 255 0 18 37
0 16 29 18 19 20 17 25 26 27
28 21 22 23 24 18 19 20 17
0
0 0 13040 0
7 74LS273
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
7931 0 0
0
0
7 Buffer~
58 161 158 0 2 22
0 30 29
0
0 0 624 270
4 4050
-14 -19 14 -11
3 U1A
13 -5 34 3
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 1 0
1 U
9325 0 0
0
0
10 Ascii Key~
169 182 99 0 11 12
0 28 27 26 25 45 46 47 30 0
0 56
0
0 0 4656 0
0
4 KBD1
-14 -34 14 -26
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
8903 0 0
0
0
9 CA 7-Seg~
184 1050 138 0 18 19
10 37 36 35 34 33 32 31 48 38
0 2 0 0 2 0 0 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3834 0 0
0
0
2 +V
167 1050 34 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3363 0 0
0
0
6 74LS47
187 1035 219 0 14 29
0 15 14 13 12 49 50 31 32 33
34 35 36 37 51
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U2
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
7668 0 0
0
0
9 Resistor~
219 1050 72 0 4 5
0 38 3 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4718 0 0
0
0
49
0 1 4 0 0 4224 0 0 6 3 0 4
790 445
790 156
945 156
945 148
3 7 4 0 0 0 0 2 7 0 0 3
722 619
722 454
843 454
3 6 4 0 0 0 0 2 7 0 0 3
722 619
722 445
843 445
3 1 5 0 0 4224 0 3 2 0 0 3
665 580
665 613
677 613
14 2 6 0 0 4224 0 9 2 0 0 3
608 391
608 625
677 625
3 2 7 0 0 4224 0 4 3 0 0 4
650 507
650 527
659 527
659 535
10 1 8 0 0 12288 0 9 3 0 0 6
662 391
662 451
677 451
677 527
671 527
671 535
11 1 9 0 0 4096 0 9 4 0 0 4
653 391
653 447
656 447
656 462
12 2 10 0 0 4096 0 9 4 0 0 2
644 391
644 462
9 1 2 0 0 8192 0 7 5 0 0 3
843 481
832 481
832 495
8 1 2 0 0 8192 0 7 5 0 0 3
843 463
832 463
832 495
5 1 2 0 0 8320 0 7 5 0 0 3
843 436
832 436
832 495
13 4 11 0 0 8320 0 9 7 0 0 3
635 391
635 427
843 427
12 3 10 0 0 8320 0 9 7 0 0 3
644 391
644 418
843 418
11 2 9 0 0 8320 0 9 7 0 0 3
653 391
653 409
843 409
10 1 8 0 0 8320 0 9 7 0 0 3
662 391
662 400
843 400
13 4 12 0 0 8320 0 7 15 0 0 3
907 454
1049 454
1049 256
12 3 13 0 0 8320 0 7 15 0 0 3
907 445
1058 445
1058 256
11 2 14 0 0 8320 0 7 15 0 0 3
907 436
1067 436
1067 256
10 1 15 0 0 8320 0 7 15 0 0 3
907 427
1076 427
1076 256
1 1 16 0 0 8320 0 1 10 0 0 4
312 203
325 203
325 219
333 219
1 9 2 0 0 0 0 8 9 0 0 4
566 332
566 319
608 319
608 327
18 6 17 0 0 12288 0 10 10 0 0 6
403 300
407 300
407 315
325 315
325 264
339 264
15 3 18 0 0 12288 0 10 10 0 0 6
403 273
407 273
407 199
325 199
325 237
339 237
16 4 19 0 0 8192 0 10 10 0 0 6
403 282
407 282
407 199
325 199
325 246
339 246
17 5 20 0 0 8192 0 10 10 0 0 6
403 291
407 291
407 199
325 199
325 255
339 255
11 1 21 0 0 4224 0 10 9 0 0 3
403 237
689 237
689 327
12 2 22 0 0 4224 0 10 9 0 0 3
403 246
680 246
680 327
13 3 23 0 0 4224 0 10 9 0 0 3
403 255
671 255
671 327
14 4 24 0 0 4224 0 10 9 0 0 3
403 264
662 264
662 327
15 5 18 0 0 4224 0 10 9 0 0 3
403 273
653 273
653 327
16 6 19 0 0 4224 0 10 9 0 0 3
403 282
644 282
644 327
17 7 20 0 0 4224 0 10 9 0 0 3
403 291
635 291
635 327
18 8 17 0 0 4224 0 10 9 0 0 3
403 300
626 300
626 327
4 7 25 0 0 8320 0 12 10 0 0 3
185 123
185 273
339 273
3 8 26 0 0 4224 0 12 10 0 0 3
191 123
191 282
339 282
2 9 27 0 0 4224 0 12 10 0 0 3
197 123
197 291
339 291
1 10 28 0 0 4224 0 12 10 0 0 3
203 123
203 300
339 300
2 2 29 0 0 8320 0 11 10 0 0 3
161 173
161 228
339 228
8 1 30 0 0 4224 0 12 11 0 0 2
161 123
161 143
7 7 31 0 0 8320 0 15 13 0 0 4
1076 186
1076 182
1065 182
1065 174
8 6 32 0 0 8320 0 15 13 0 0 4
1067 186
1067 182
1059 182
1059 174
9 5 33 0 0 12416 0 15 13 0 0 4
1058 186
1058 182
1053 182
1053 174
10 4 34 0 0 12416 0 15 13 0 0 4
1049 186
1049 182
1047 182
1047 174
11 3 35 0 0 12416 0 15 13 0 0 4
1040 186
1040 182
1041 182
1041 174
12 2 36 0 0 12416 0 15 13 0 0 4
1031 186
1031 182
1035 182
1035 174
13 1 37 0 0 12416 0 15 13 0 0 4
1022 186
1022 182
1029 182
1029 174
1 2 3 0 0 4224 0 14 16 0 0 2
1050 43
1050 54
1 9 38 0 0 4224 0 16 13 0 0 2
1050 90
1050 102
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
