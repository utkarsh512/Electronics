CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 7 100 9
38 96 1498 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 96 1498 799
143654930 0
0
6 Title:
5 Name:
0
0
0
39
13 Logic Switch~
5 607 454 0 10 11
0 29 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-32 6 -18 14
3 V11
-35 -5 -14 3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 252 172 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-32 6 -18 14
3 V10
-35 -5 -14 3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 252 202 0 1 11
0 27
0
0 0 21360 0
2 0V
-32 6 -18 14
2 V9
-32 -5 -18 3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 252 236 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-32 6 -18 14
2 V8
-32 -5 -18 3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 253 269 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-32 6 -18 14
2 V7
-32 -5 -18 3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 708 126 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
22 0 36 8
2 V6
22 -9 36 -1
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 708 99 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
22 0 36 8
2 V5
22 -9 36 -1
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 706 69 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
22 0 36 8
2 V4
22 -9 36 -1
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3747 0 0
0
0
13 Logic Switch~
5 705 42 0 1 11
0 21
0
0 0 21360 512
2 0V
19 -5 33 3
2 V3
19 -16 33 -8
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3549 0 0
0
0
13 Logic Switch~
5 72 27 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7931 0 0
0
0
13 Logic Switch~
5 517 21 0 1 11
0 32
0
0 0 21360 512
2 0V
-7 21 7 29
2 V1
-7 10 7 18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9325 0 0
0
0
14 Logic Display~
6 436 202 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8903 0 0
0
0
14 Logic Display~
6 418 202 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3834 0 0
0
0
14 Logic Display~
6 401 202 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3363 0 0
0
0
14 Logic Display~
6 384 202 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7668 0 0
0
0
14 Logic Display~
6 490 205 0 1 2
10 3
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L10
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4718 0 0
0
0
14 Logic Display~
6 212 68 0 1 2
10 8
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L9
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3874 0 0
0
0
14 Logic Display~
6 310 373 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6671 0 0
0
0
14 Logic Display~
6 264 457 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3789 0 0
0
0
14 Logic Display~
6 285 460 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4871 0 0
0
0
14 Logic Display~
6 306 460 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3750 0 0
0
0
14 Logic Display~
6 327 459 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8778 0 0
0
0
14 Logic Display~
6 350 460 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
538 0 0
0
0
14 Logic Display~
6 370 461 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6843 0 0
0
0
14 Logic Display~
6 391 462 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3136 0 0
0
0
14 Logic Display~
6 410 460 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5950 0 0
0
0
9 2-In AND~
219 534 207 0 3 22
0 3 21 17
0
0 0 624 782
6 74LS08
-21 -24 21 -16
3 U6D
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 2 0
1 U
5670 0 0
0
0
9 2-In AND~
219 571 207 0 3 22
0 3 22 18
0
0 0 624 782
6 74LS08
-21 -24 21 -16
3 U6C
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 2 0
1 U
6828 0 0
0
0
9 2-In AND~
219 611 208 0 3 22
0 3 23 19
0
0 0 624 782
6 74LS08
-21 -24 21 -16
3 U6B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 2 0
1 U
6735 0 0
0
0
9 2-In AND~
219 654 209 0 3 22
0 3 24 20
0
0 0 624 782
6 74LS08
-21 -24 21 -16
3 U6A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 1803067004
65 0 0 0 4 1 2 0
1 U
8365 0 0
0
0
7 Ground~
168 396 151 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4132 0 0
0
0
9 Inverter~
13 133 237 0 2 22
0 30 7
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U5C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 3 1 0
1 U
4551 0 0
0
0
9 Inverter~
13 133 183 0 2 22
0 31 30
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U5B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 1 0
1 U
3635 0 0
0
0
9 Inverter~
13 134 128 0 2 22
0 8 31
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U5A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 1 0
1 U
3973 0 0
0
0
6 74LS95
110 459 131 0 12 25
0 32 8 8 25 26 27 28 2 3
4 5 6
0
0 0 13040 270
6 74LS95
-21 -51 21 -43
2 U4
45 0 59 8
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 6 9 8 5 4 3 2 1 10
11 12 13 6 9 8 5 4 3 2
1 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
3851 0 0
0
0
7 Ground~
168 893 274 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8383 0 0
0
0
7 74LS273
150 732 454 0 18 37
0 29 7 34 35 36 37 38 39 40
41 9 10 11 12 13 14 15 16
0
0 0 13040 782
7 74LS273
-24 -60 25 -52
2 U3
54 0 68 8
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
9334 0 0
0
0
6 74LS83
105 650 296 0 14 29
0 9 10 11 12 17 18 19 20 33
35 36 37 38 34
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
2 U2
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
7471 0 0
0
0
6 74LS83
105 816 297 0 14 29
0 13 14 15 16 2 2 2 2 2
39 40 41 42 33
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
2 U1
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3334 0 0
0
0
62
9 1 3 0 0 4096 0 35 12 0 0 4
449 168
449 228
436 228
436 220
10 1 4 0 0 8320 0 35 13 0 0 6
440 168
440 187
371 187
371 228
418 228
418 220
11 1 5 0 0 8320 0 35 14 0 0 6
431 168
431 187
371 187
371 228
401 228
401 220
12 1 6 0 0 8320 0 35 15 0 0 6
422 168
422 187
371 187
371 228
384 228
384 220
1 0 7 0 0 4096 0 18 0 0 42 2
310 391
310 413
1 0 3 0 0 0 0 16 0 0 31 4
490 191
490 184
491 184
491 179
1 0 8 0 0 4096 0 17 0 0 46 2
212 54
212 27
11 1 9 0 0 8320 0 37 19 0 0 4
709 491
709 637
264 637
264 475
12 1 10 0 0 8320 0 37 20 0 0 4
718 491
718 629
285 629
285 478
13 1 11 0 0 8320 0 37 21 0 0 4
727 491
727 621
306 621
306 478
14 1 12 0 0 8320 0 37 22 0 0 4
736 491
736 614
327 614
327 477
15 1 13 0 0 8320 0 37 23 0 0 4
745 491
745 607
350 607
350 478
16 1 14 0 0 8320 0 37 24 0 0 4
754 491
754 600
370 600
370 479
17 1 15 0 0 8320 0 37 25 0 0 4
763 491
763 594
391 594
391 480
18 1 16 0 0 8320 0 37 26 0 0 4
772 491
772 587
410 587
410 478
15 1 13 0 0 12416 0 37 39 0 0 6
745 491
745 557
1068 557
1068 134
778 134
778 267
16 2 14 0 0 12416 0 37 39 0 0 6
754 491
754 537
1054 537
1054 140
787 140
787 267
17 3 15 0 0 0 0 37 39 0 0 6
763 491
763 519
1039 519
1039 148
796 148
796 267
18 4 16 0 0 0 0 37 39 0 0 6
772 491
772 495
1024 495
1024 159
805 159
805 267
14 4 12 0 0 0 0 37 38 0 0 6
736 491
736 558
433 558
433 250
639 250
639 266
13 3 11 0 0 0 0 37 38 0 0 6
727 491
727 537
480 537
480 253
630 253
630 266
12 2 10 0 0 0 0 37 38 0 0 6
718 491
718 520
524 520
524 256
621 256
621 266
11 1 9 0 0 0 0 37 38 0 0 8
709 491
709 495
550 495
550 334
551 334
551 260
612 260
612 266
3 5 17 0 0 8320 0 27 38 0 0 4
532 230
532 247
648 247
648 266
3 6 18 0 0 8320 0 28 38 0 0 4
569 230
569 244
657 244
657 266
3 7 19 0 0 8320 0 29 38 0 0 4
609 231
609 241
666 241
666 266
3 8 20 0 0 12416 0 30 38 0 0 4
652 232
652 238
675 238
675 266
1 0 3 0 0 0 0 27 0 0 31 2
523 185
523 179
1 0 3 0 0 0 0 28 0 0 31 2
560 185
560 179
1 0 3 0 0 0 0 29 0 0 31 3
600 186
600 179
601 179
9 1 3 0 0 8320 0 35 30 0 0 4
449 168
449 179
643 179
643 187
1 2 21 0 0 4224 0 9 27 0 0 3
693 42
541 42
541 185
1 2 22 0 0 4224 0 8 28 0 0 3
694 69
578 69
578 185
1 2 23 0 0 8320 0 7 29 0 0 3
696 99
618 99
618 186
1 2 24 0 0 8320 0 6 30 0 0 3
696 126
661 126
661 187
8 1 2 0 0 12288 0 35 31 0 0 4
422 104
422 98
396 98
396 145
1 4 25 0 0 8320 0 5 35 0 0 5
265 269
365 269
365 90
458 90
458 104
1 5 26 0 0 8320 0 4 35 0 0 5
264 236
343 236
343 67
449 67
449 104
1 6 27 0 0 8320 0 3 35 0 0 5
264 202
323 202
323 53
440 53
440 104
1 7 28 0 0 8320 0 2 35 0 0 5
264 172
305 172
305 37
431 37
431 104
1 1 29 0 0 12416 0 1 37 0 0 5
619 454
633 454
633 422
691 422
691 421
2 2 7 0 0 8320 0 32 37 0 0 4
136 255
136 413
700 413
700 427
2 1 30 0 0 4224 0 33 32 0 0 2
136 201
136 219
2 1 31 0 0 4224 0 34 33 0 0 4
137 146
137 157
136 157
136 165
1 1 8 0 0 4096 0 34 10 0 0 3
137 110
137 27
84 27
1 0 8 0 0 4224 0 10 0 0 47 3
84 27
471 27
471 98
3 2 8 0 0 0 0 35 35 0 0 2
467 98
476 98
1 1 32 0 0 8320 0 11 35 0 0 3
505 21
485 21
485 104
5 1 2 0 0 12416 0 39 36 0 0 4
814 267
814 188
893 188
893 268
6 1 2 0 0 0 0 39 36 0 0 4
823 267
823 208
893 208
893 268
7 1 2 0 0 0 0 39 36 0 0 4
832 267
832 222
893 222
893 268
8 1 2 0 0 0 0 39 36 0 0 4
841 267
841 235
893 235
893 268
9 1 2 0 0 0 0 39 36 0 0 4
859 267
859 260
893 260
893 268
9 14 33 0 0 8320 0 38 39 0 0 6
693 266
693 180
960 180
960 339
859 339
859 331
3 14 34 0 0 4224 0 37 38 0 0 4
709 427
709 338
693 338
693 330
4 10 35 0 0 8320 0 37 38 0 0 4
718 427
718 399
639 399
639 330
5 11 36 0 0 8320 0 37 38 0 0 4
727 427
727 381
648 381
648 330
6 12 37 0 0 8320 0 37 38 0 0 4
736 427
736 362
657 362
657 330
7 13 38 0 0 8320 0 37 38 0 0 4
745 427
745 350
666 350
666 330
8 10 39 0 0 12416 0 37 39 0 0 4
754 427
754 394
805 394
805 331
9 11 40 0 0 12416 0 37 39 0 0 4
763 427
763 404
814 404
814 331
12 10 41 0 0 4224 0 39 37 0 0 4
823 331
823 413
772 413
772 427
11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
1180 27 1260 51
1190 35 1262 51
9 18EC30048
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
1181 13 1293 37
1191 21 1295 37
13 UTKARSH PATEL
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
1133 199 1317 223
1143 207 1319 223
22 5. Read o/p from lamps
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
1135 173 1303 197
1145 181 1305 197
20 4. Apply CLK 4 times
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
1136 142 1248 166
1146 150 1250 166
13 3. Reset MODE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
1137 118 1321 142
1147 126 1323 142
22 2. Set MODE, apply CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
1138 95 1298 119
1148 103 1300 119
19 1. Reset and set MR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1138 53 1194 77
1148 61 1196 77
6 Steps:
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
563 463 587 487
573 471 589 487
2 MR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
535 5 575 29
545 13 577 29
4 MODE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
35 38 83 62
45 46 85 62
5 CLOCK
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
