CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
70 0 5 130 9
38 96 1497 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 96 1497 799
143654930 0
0
6 Title:
5 Name:
0
0
0
18
11 2-Input OR~
1 442 375 0 3 22
0 11 10 7
0
0 0 880 180
6 74LS32
-9 -25 33 -17
3 U7A
1 -35 22 -27
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 515768069
65 0 0 0 4 1 5 0
1 U
8953 0 0
0
0
12 2-Input AND~
0 509 368 0 3 22
0 6 12 10
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U6B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 431816451
65 0 0 0 4 2 3 0
1 U
4441 0 0
0
0
11 3-Input OR~
86 505 332 0 4 22
0 11 13 14 9
0
0 0 624 180
4 4075
-14 -28 14 -20
3 U3A
1 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 3 5 6 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 4 0
1 U
3618 0 0
0
0
12 2-Input AND~
0 912 393 0 3 22
0 15 16 6
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U6A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 3 0
1 U
6153 0 0
0
0
12 2-Input AND~
0 847 391 0 3 22
0 17 15 8
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U4D
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 1 0
1 U
5394 0 0
0
0
12 2-Input AND~
0 781 392 0 3 22
0 17 18 11
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U4C
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 1 0
1 U
7734 0 0
0
0
12 2-Input AND~
0 711 392 0 3 22
0 4 18 13
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U4B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 314375944
65 0 0 0 4 2 1 0
1 U
9914 0 0
0
0
13 2-Input NAND~
2 695 308 0 3 22
0 12 12 18
0
0 0 880 270
6 74LS00
20 -2 62 6
3 U5C
30 -12 51 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 2 0
1 U
3747 0 0
0
0
13 2-Input NAND~
2 736 308 0 3 22
0 17 17 16
0
0 0 880 270
6 74LS00
20 -2 62 6
3 U5B
30 -12 51 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 2 0
1 U
3549 0 0
0
0
13 2-Input NAND~
2 776 308 0 3 22
0 4 4 15
0
0 0 880 270
6 74LS00
20 -2 62 6
3 U5A
30 -12 51 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 314375944
65 0 0 0 4 1 2 0
1 U
7931 0 0
0
0
12 2-Input AND~
0 862 261 0 3 22
0 4 17 14
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U4A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 431816451
65 0 0 0 4 1 1 0
1 U
9325 0 0
0
0
7 Pulser~
4 823 95 0 10 12
0 27 28 5 29 0 0 5 5 2
7
0
0 0 4656 512
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
8903 0 0
0
0
7 Ground~
168 707 115 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3834 0 0
0
0
6 74LS93
109 756 157 0 8 17
0 2 2 5 4 30 12 17 4
0
0 0 13040 782
6 74LS93
-21 -35 21 -27
2 U2
28 0 42 8
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 512 1 0 0 0
1 U
3363 0 0
0
0
6 74LS47
187 389 262 0 14 29
0 9 8 7 6 31 32 19 20 21
22 23 24 25 33
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U1
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
7668 0 0
0
0
2 +V
167 404 77 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4718 0 0
0
0
9 CA 7-Seg~
184 404 181 0 18 19
10 25 24 23 22 21 20 19 34 26
2 0 0 2 2 2 2 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3874 0 0
0
0
9 Resistor~
219 404 115 0 4 5
0 26 3 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6671 0 0
0
0
40
8 4 4 0 0 12288 0 14 14 0 0 6
770 193
770 197
785 197
785 115
770 115
770 123
3 3 5 0 0 8320 0 14 12 0 0 3
761 123
761 86
799 86
4 3 6 0 0 8320 0 15 4 0 0 4
403 299
403 424
910 424
910 416
3 3 7 0 0 4224 0 15 1 0 0 3
412 299
412 375
415 375
2 3 8 0 0 8320 0 15 5 0 0 4
421 299
421 422
845 422
845 414
1 4 9 0 0 8320 0 15 3 0 0 3
430 299
430 332
478 332
2 3 10 0 0 4240 0 1 2 0 0 4
460 369
478 369
478 368
482 368
3 1 11 0 0 8320 0 6 1 0 0 5
779 415
779 419
482 419
482 381
460 381
1 3 6 0 0 0 0 2 4 0 0 5
527 374
690 374
690 424
910 424
910 416
6 2 12 0 0 8320 0 14 2 0 0 5
752 193
752 279
543 279
543 362
527 362
3 1 11 0 0 0 0 6 3 0 0 5
779 415
779 419
546 419
546 341
524 341
3 2 13 0 0 8320 0 7 3 0 0 5
709 415
709 419
546 419
546 332
523 332
3 3 14 0 0 8320 0 11 3 0 0 5
860 284
860 339
546 339
546 323
524 323
3 1 15 0 0 8320 0 10 4 0 0 4
777 334
777 363
916 363
916 371
3 2 16 0 0 8320 0 9 4 0 0 4
737 334
737 363
904 363
904 371
3 2 15 0 0 0 0 10 5 0 0 4
777 334
777 361
839 361
839 369
7 1 17 0 0 4096 0 14 5 0 0 6
761 193
761 279
841 279
841 289
851 289
851 369
7 1 17 0 0 0 0 14 6 0 0 6
761 193
761 279
797 279
797 362
785 362
785 370
3 2 18 0 0 12416 0 8 6 0 0 5
696 334
703 334
703 348
773 348
773 370
8 1 4 0 0 16384 0 14 7 0 0 5
770 193
766 193
766 279
715 279
715 370
3 2 18 0 0 0 0 8 7 0 0 4
696 334
696 362
703 362
703 370
8 0 4 0 0 0 0 14 0 0 25 3
770 193
770 193
771 275
7 0 17 0 0 0 0 14 0 0 26 4
761 193
761 270
740 270
740 275
6 0 12 0 0 0 0 14 0 0 27 4
752 193
752 208
695 208
695 275
2 1 4 0 0 0 0 10 10 0 0 4
771 283
771 275
783 275
783 283
2 1 17 0 0 0 0 9 9 0 0 4
731 283
731 275
743 275
743 283
2 1 12 0 0 0 0 8 8 0 0 4
690 283
690 275
702 275
702 283
7 2 17 0 0 8320 0 14 11 0 0 4
761 193
761 207
854 207
854 239
8 1 4 0 0 8320 0 14 11 0 0 4
770 193
770 199
866 199
866 239
0 1 2 0 0 4224 0 0 13 31 0 4
747 129
747 85
707 85
707 109
1 2 2 0 0 0 0 14 14 0 0 2
743 129
752 129
7 7 19 0 0 8320 0 15 17 0 0 4
430 229
430 225
419 225
419 217
8 6 20 0 0 8320 0 15 17 0 0 4
421 229
421 225
413 225
413 217
9 5 21 0 0 12416 0 15 17 0 0 4
412 229
412 225
407 225
407 217
10 4 22 0 0 12416 0 15 17 0 0 4
403 229
403 225
401 225
401 217
11 3 23 0 0 12416 0 15 17 0 0 4
394 229
394 225
395 225
395 217
12 2 24 0 0 12416 0 15 17 0 0 4
385 229
385 225
389 225
389 217
13 1 25 0 0 12416 0 15 17 0 0 4
376 229
376 225
383 225
383 217
1 2 3 0 0 4224 0 16 18 0 0 2
404 86
404 97
1 9 26 0 0 4224 0 18 17 0 0 2
404 133
404 145
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
899 378 923 402
907 384 923 400
2 ba
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
824 383 848 407
832 389 848 405
2 Ba
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
748 383 772 407
755 389 771 405
2 cB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
666 375 690 399
674 381 690 397
2 cA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
791 319 815 343
798 325 814 341
2 A_
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
712 319 736 343
720 325 736 341
2 B_
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
654 313 678 337
662 319 678 335
2 c_
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
878 275 902 299
885 281 901 297
2 BA
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
